

    module uriscv_csr_SUPPORT_CSR1_SUPPORT_MCYCLE1_SUPPORT_MTIMECMP0_SUPPORT_MSCRATCH0_SUPPORT_MIP_MIE0_SUPPORT_MTVEC0_SUPPORT_MTVAL0_SUPPORT_MULDIV1 ( 
        clk_i, rst_i, intr_i, isr_vector_i, cpu_id_i, valid_i, pc_i, opcode_i, 
        rs1_val_i, rs2_val_i, csr_rdata_o, excpn_invalid_inst_i, 
        excpn_lsu_align_i, mem_addr_i, csr_mepc_o, exception_o, 
        exception_type_o, exception_pc_o );
  input [31:0] isr_vector_i;
  input [31:0] cpu_id_i;
  input [31:0] pc_i;
  input [31:0] opcode_i;
  input [31:0] rs1_val_i;
  input [31:0] rs2_val_i;
  output [31:0] csr_rdata_o;
  input [31:0] mem_addr_i;
  output [31:0] csr_mepc_o;
  output [5:0] exception_type_o;
  output [31:0] exception_pc_o;
  input clk_i, rst_i, intr_i, valid_i, excpn_invalid_inst_i, excpn_lsu_align_i;
  output exception_o;
  wire   csr_mcause_r_31_, N818, N819, N820, N821, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n74, n75, n118, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n1, n2, n3, n20, n21, n79,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450;
  wire   [31:0] csr_mcause_q;
  wire   [31:0] csr_sr_q;
  wire   [31:0] csr_mcycle_q;
  wire   [31:4] csr_mcycle_r;

  DFF_X1 csr_mcause_q_reg_3_ ( .D(N821), .CK(clk_i), .Q(csr_mcause_q[3]), .QN(
        n97) );
  DFF_X1 csr_mcause_q_reg_1_ ( .D(N819), .CK(clk_i), .Q(csr_mcause_q[1]), .QN(
        n105) );
  DFF_X1 csr_mcause_q_reg_0_ ( .D(N818), .CK(clk_i), .Q(csr_mcause_q[0]), .QN(
        n103) );
  SDFF_X1 csr_mcause_q_reg_31_ ( .D(1'b0), .SI(n118), .SE(csr_mcause_r_31_), 
        .CK(clk_i), .Q(csr_mcause_q[31]), .QN(n104) );
  DFF_X1 csr_mcause_q_reg_2_ ( .D(N820), .CK(clk_i), .Q(csr_mcause_q[2]), .QN(
        n96) );
  DFF_X1 csr_mepc_q_reg_1_ ( .D(n618), .CK(clk_i), .Q(csr_mepc_o[1]), .QN(n75)
         );
  DFF_X1 csr_mepc_q_reg_2_ ( .D(n617), .CK(clk_i), .Q(csr_mepc_o[2]), .QN(n74)
         );
  DFF_X1 csr_mepc_q_reg_5_ ( .D(n614), .CK(clk_i), .Q(csr_mepc_o[5]), .QN(n71)
         );
  DFF_X1 csr_mepc_q_reg_6_ ( .D(n613), .CK(clk_i), .Q(csr_mepc_o[6]), .QN(n70)
         );
  DFF_X1 csr_mepc_q_reg_7_ ( .D(n612), .CK(clk_i), .Q(csr_mepc_o[7]), .QN(n69)
         );
  DFF_X1 csr_mepc_q_reg_8_ ( .D(n611), .CK(clk_i), .Q(csr_mepc_o[8]), .QN(n68)
         );
  DFF_X1 csr_mepc_q_reg_9_ ( .D(n610), .CK(clk_i), .Q(csr_mepc_o[9]), .QN(n67)
         );
  DFF_X1 csr_mepc_q_reg_10_ ( .D(n609), .CK(clk_i), .Q(csr_mepc_o[10]), .QN(
        n66) );
  DFF_X1 csr_mepc_q_reg_11_ ( .D(n608), .CK(clk_i), .Q(csr_mepc_o[11]), .QN(
        n65) );
  DFF_X1 csr_mepc_q_reg_12_ ( .D(n607), .CK(clk_i), .Q(csr_mepc_o[12]), .QN(
        n64) );
  DFF_X1 csr_mepc_q_reg_13_ ( .D(n606), .CK(clk_i), .Q(csr_mepc_o[13]), .QN(
        n63) );
  DFF_X1 csr_mepc_q_reg_14_ ( .D(n605), .CK(clk_i), .Q(csr_mepc_o[14]), .QN(
        n62) );
  DFF_X1 csr_mepc_q_reg_15_ ( .D(n604), .CK(clk_i), .Q(csr_mepc_o[15]), .QN(
        n61) );
  DFF_X1 csr_mepc_q_reg_16_ ( .D(n603), .CK(clk_i), .Q(csr_mepc_o[16]), .QN(
        n60) );
  DFF_X1 csr_mepc_q_reg_17_ ( .D(n602), .CK(clk_i), .Q(csr_mepc_o[17]), .QN(
        n59) );
  DFF_X1 csr_mepc_q_reg_18_ ( .D(n601), .CK(clk_i), .Q(csr_mepc_o[18]), .QN(
        n58) );
  DFF_X1 csr_mepc_q_reg_19_ ( .D(n600), .CK(clk_i), .Q(csr_mepc_o[19]), .QN(
        n57) );
  DFF_X1 csr_mepc_q_reg_20_ ( .D(n599), .CK(clk_i), .Q(csr_mepc_o[20]), .QN(
        n56) );
  DFF_X1 csr_mepc_q_reg_21_ ( .D(n598), .CK(clk_i), .Q(csr_mepc_o[21]), .QN(
        n55) );
  DFF_X1 csr_mepc_q_reg_22_ ( .D(n597), .CK(clk_i), .Q(csr_mepc_o[22]), .QN(
        n54) );
  DFF_X1 csr_mepc_q_reg_23_ ( .D(n596), .CK(clk_i), .Q(csr_mepc_o[23]), .QN(
        n53) );
  DFF_X1 csr_mepc_q_reg_24_ ( .D(n595), .CK(clk_i), .Q(csr_mepc_o[24]), .QN(
        n52) );
  DFF_X1 csr_mepc_q_reg_25_ ( .D(n594), .CK(clk_i), .Q(csr_mepc_o[25]), .QN(
        n51) );
  DFF_X1 csr_mepc_q_reg_26_ ( .D(n593), .CK(clk_i), .Q(csr_mepc_o[26]), .QN(
        n50) );
  DFF_X1 csr_mepc_q_reg_27_ ( .D(n592), .CK(clk_i), .Q(csr_mepc_o[27]), .QN(
        n49) );
  DFF_X1 csr_mepc_q_reg_28_ ( .D(n591), .CK(clk_i), .Q(csr_mepc_o[28]), .QN(
        n48) );
  DFF_X1 csr_mepc_q_reg_29_ ( .D(n590), .CK(clk_i), .Q(csr_mepc_o[29]), .QN(
        n47) );
  DFF_X1 csr_mepc_q_reg_30_ ( .D(n589), .CK(clk_i), .Q(csr_mepc_o[30]), .QN(
        n46) );
  DFF_X1 csr_mepc_q_reg_31_ ( .D(n588), .CK(clk_i), .Q(csr_mepc_o[31]), .QN(
        n45) );
  DFF_X1 csr_sr_q_reg_7_ ( .D(n584), .CK(clk_i), .Q(csr_sr_q[7]), .QN(n106) );
  SDFF_X1 csr_mcycle_q_reg_29_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[29]), 
        .CK(clk_i), .Q(csr_mcycle_q[29]), .QN(n99) );
  SDFF_X1 csr_mcycle_q_reg_27_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[27]), 
        .CK(clk_i), .Q(csr_mcycle_q[27]), .QN(n100) );
  SDFF_X1 csr_mcycle_q_reg_25_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[25]), 
        .CK(clk_i), .Q(csr_mcycle_q[25]), .QN(n101) );
  SDFF_X1 csr_mcycle_q_reg_23_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[23]), 
        .CK(clk_i), .Q(csr_mcycle_q[23]), .QN(n102) );
  SDFF_X1 csr_mcycle_q_reg_21_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[21]), 
        .CK(clk_i), .Q(csr_mcycle_q[21]), .QN(n87) );
  SDFF_X1 csr_mcycle_q_reg_19_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[19]), 
        .CK(clk_i), .Q(csr_mcycle_q[19]), .QN(n88) );
  SDFF_X1 csr_mcycle_q_reg_17_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[17]), 
        .CK(clk_i), .Q(csr_mcycle_q[17]), .QN(n89) );
  SDFF_X1 csr_mcycle_q_reg_15_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[15]), 
        .CK(clk_i), .Q(csr_mcycle_q[15]), .QN(n90) );
  SDFF_X1 csr_mcycle_q_reg_13_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[13]), 
        .CK(clk_i), .Q(csr_mcycle_q[13]), .QN(n91) );
  SDFF_X1 csr_mcycle_q_reg_11_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[11]), 
        .CK(clk_i), .Q(csr_mcycle_q[11]), .QN(n92) );
  SDFF_X1 csr_mcycle_q_reg_9_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[9]), 
        .CK(clk_i), .Q(csr_mcycle_q[9]), .QN(n93) );
  SDFF_X1 csr_mcycle_q_reg_7_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[7]), 
        .CK(clk_i), .Q(csr_mcycle_q[7]), .QN(n94) );
  SDFF_X1 csr_mcycle_q_reg_5_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[5]), 
        .CK(clk_i), .Q(csr_mcycle_q[5]), .QN(n95) );
  SDFF_X1 csr_mcycle_q_reg_0_ ( .D(1'b0), .SI(n118), .SE(n85), .CK(clk_i), .Q(
        csr_mcycle_q[0]), .QN(n85) );
  DFF_X1 csr_mcycle_q_reg_3_ ( .D(n21), .CK(clk_i), .QN(n86) );
  DFF_X1 csr_mcycle_q_reg_1_ ( .D(n20), .CK(clk_i), .Q(csr_mcycle_q[1]), .QN(
        n98) );
  SDFF_X1 csr_mcycle_q_reg_2_ ( .D(n118), .SI(1'b0), .SE(n142), .CK(clk_i), 
        .Q(csr_mcycle_q[2]) );
  SDFF_X1 csr_mcycle_q_reg_4_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[4]), 
        .CK(clk_i), .Q(csr_mcycle_q[4]) );
  SDFF_X1 csr_mcycle_q_reg_6_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[6]), 
        .CK(clk_i), .Q(csr_mcycle_q[6]) );
  SDFF_X1 csr_mcycle_q_reg_8_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[8]), 
        .CK(clk_i), .Q(csr_mcycle_q[8]) );
  SDFF_X1 csr_mcycle_q_reg_10_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[10]), 
        .CK(clk_i), .Q(csr_mcycle_q[10]) );
  SDFF_X1 csr_mcycle_q_reg_12_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[12]), 
        .CK(clk_i), .Q(csr_mcycle_q[12]) );
  SDFF_X1 csr_mcycle_q_reg_14_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[14]), 
        .CK(clk_i), .Q(csr_mcycle_q[14]) );
  SDFF_X1 csr_mcycle_q_reg_16_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[16]), 
        .CK(clk_i), .Q(csr_mcycle_q[16]) );
  SDFF_X1 csr_mcycle_q_reg_18_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[18]), 
        .CK(clk_i), .Q(csr_mcycle_q[18]) );
  SDFF_X1 csr_mcycle_q_reg_20_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[20]), 
        .CK(clk_i), .Q(csr_mcycle_q[20]) );
  SDFF_X1 csr_mcycle_q_reg_22_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[22]), 
        .CK(clk_i), .Q(csr_mcycle_q[22]) );
  SDFF_X1 csr_mcycle_q_reg_24_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[24]), 
        .CK(clk_i), .Q(csr_mcycle_q[24]) );
  SDFF_X1 csr_mcycle_q_reg_26_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[26]), 
        .CK(clk_i), .Q(csr_mcycle_q[26]) );
  SDFF_X1 csr_mcycle_q_reg_28_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[28]), 
        .CK(clk_i), .Q(csr_mcycle_q[28]) );
  SDFF_X1 csr_mcycle_q_reg_30_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[30]), 
        .CK(clk_i), .Q(csr_mcycle_q[30]) );
  SDFF_X1 csr_mcycle_q_reg_31_ ( .D(1'b0), .SI(n118), .SE(csr_mcycle_r[31]), 
        .CK(clk_i), .Q(csr_mcycle_q[31]) );
  DFF_X1 csr_sr_q_reg_3_ ( .D(n622), .CK(clk_i), .Q(csr_sr_q[3]) );
  DFF_X1 csr_sr_q_reg_1_ ( .D(n620), .CK(clk_i), .Q(csr_sr_q[1]) );
  DFF_X1 csr_sr_q_reg_0_ ( .D(n623), .CK(clk_i), .Q(csr_sr_q[0]) );
  DFF_X1 csr_sr_q_reg_2_ ( .D(n621), .CK(clk_i), .Q(csr_sr_q[2]) );
  DFF_X1 csr_sr_q_reg_4_ ( .D(n587), .CK(clk_i), .Q(csr_sr_q[4]) );
  DFF_X1 csr_sr_q_reg_31_ ( .D(n560), .CK(clk_i), .Q(csr_sr_q[31]) );
  DFF_X1 csr_mepc_q_reg_0_ ( .D(n619), .CK(clk_i), .Q(csr_mepc_o[0]) );
  DFF_X1 csr_mepc_q_reg_3_ ( .D(n616), .CK(clk_i), .Q(csr_mepc_o[3]) );
  DFF_X1 csr_mepc_q_reg_4_ ( .D(n615), .CK(clk_i), .Q(csr_mepc_o[4]) );
  DFF_X1 csr_sr_q_reg_12_ ( .D(n579), .CK(clk_i), .Q(csr_sr_q[12]) );
  DFF_X1 csr_sr_q_reg_11_ ( .D(n580), .CK(clk_i), .Q(csr_sr_q[11]) );
  DFF_X1 csr_sr_q_reg_26_ ( .D(n565), .CK(clk_i), .Q(csr_sr_q[26]) );
  DFF_X1 csr_sr_q_reg_23_ ( .D(n568), .CK(clk_i), .Q(csr_sr_q[23]) );
  DFF_X1 csr_sr_q_reg_21_ ( .D(n570), .CK(clk_i), .Q(csr_sr_q[21]) );
  DFF_X1 csr_sr_q_reg_19_ ( .D(n572), .CK(clk_i), .Q(csr_sr_q[19]) );
  DFF_X1 csr_sr_q_reg_18_ ( .D(n573), .CK(clk_i), .Q(csr_sr_q[18]) );
  DFF_X1 csr_sr_q_reg_17_ ( .D(n574), .CK(clk_i), .Q(csr_sr_q[17]) );
  DFF_X1 csr_sr_q_reg_16_ ( .D(n575), .CK(clk_i), .Q(csr_sr_q[16]) );
  DFF_X1 csr_sr_q_reg_15_ ( .D(n576), .CK(clk_i), .Q(csr_sr_q[15]) );
  DFF_X1 csr_sr_q_reg_9_ ( .D(n582), .CK(clk_i), .Q(csr_sr_q[9]) );
  DFF_X1 csr_sr_q_reg_8_ ( .D(n583), .CK(clk_i), .Q(csr_sr_q[8]) );
  DFF_X1 csr_sr_q_reg_6_ ( .D(n585), .CK(clk_i), .Q(csr_sr_q[6]) );
  DFF_X1 csr_sr_q_reg_5_ ( .D(n586), .CK(clk_i), .Q(csr_sr_q[5]) );
  DFF_X1 csr_sr_q_reg_30_ ( .D(n561), .CK(clk_i), .Q(csr_sr_q[30]) );
  DFF_X1 csr_sr_q_reg_29_ ( .D(n562), .CK(clk_i), .Q(csr_sr_q[29]) );
  DFF_X1 csr_sr_q_reg_28_ ( .D(n563), .CK(clk_i), .Q(csr_sr_q[28]) );
  DFF_X1 csr_sr_q_reg_27_ ( .D(n564), .CK(clk_i), .Q(csr_sr_q[27]) );
  DFF_X1 csr_sr_q_reg_25_ ( .D(n566), .CK(clk_i), .Q(csr_sr_q[25]) );
  DFF_X1 csr_sr_q_reg_24_ ( .D(n567), .CK(clk_i), .Q(csr_sr_q[24]) );
  DFF_X1 csr_sr_q_reg_22_ ( .D(n569), .CK(clk_i), .Q(csr_sr_q[22]) );
  DFF_X1 csr_sr_q_reg_20_ ( .D(n571), .CK(clk_i), .Q(csr_sr_q[20]) );
  DFF_X1 csr_sr_q_reg_14_ ( .D(n577), .CK(clk_i), .Q(csr_sr_q[14]) );
  DFF_X1 csr_sr_q_reg_13_ ( .D(n578), .CK(clk_i), .Q(csr_sr_q[13]) );
  DFF_X1 csr_sr_q_reg_10_ ( .D(n581), .CK(clk_i), .Q(csr_sr_q[10]) );
  INV_X1 U3 ( .A(n118), .ZN(n1) );
  AOI211_X1 U4 ( .C1(n85), .C2(n98), .A(n143), .B(n1), .ZN(n20) );
  INV_X1 U5 ( .A(opcode_i[27]), .ZN(n2) );
  NAND3_X1 U6 ( .A1(opcode_i[26]), .A2(n208), .A3(n2), .ZN(n198) );
  INV_X1 U7 ( .A(n118), .ZN(n3) );
  AOI211_X1 U8 ( .C1(n141), .C2(n86), .A(n140), .B(n3), .ZN(n21) );
  INV_X1 U25 ( .A(n371), .ZN(n366) );
  INV_X2 U26 ( .A(n271), .ZN(n292) );
  BUF_X2 U27 ( .A(n442), .Z(n79) );
  INV_X2 U28 ( .A(n387), .ZN(n446) );
  NOR2_X1 U29 ( .A1(n146), .A2(n286), .ZN(exception_o) );
  NOR2_X1 U30 ( .A1(excpn_lsu_align_i), .A2(n83), .ZN(n146) );
  OR2_X1 U31 ( .A1(excpn_invalid_inst_i), .A2(n84), .ZN(n83) );
  INV_X2 U32 ( .A(n259), .ZN(n272) );
  BUF_X2 U33 ( .A(n273), .Z(n82) );
  AND3_X2 U34 ( .A1(n209), .A2(n208), .A3(n211), .ZN(n276) );
  AND2_X1 U35 ( .A1(intr_i), .A2(csr_sr_q[3]), .ZN(n84) );
  INV_X2 U36 ( .A(rst_i), .ZN(n118) );
  NOR4_X2 U37 ( .A1(opcode_i[22]), .A2(n157), .A3(n148), .A4(n198), .ZN(n256)
         );
  BUF_X1 U38 ( .A(n374), .Z(n112) );
  BUF_X1 U39 ( .A(n365), .Z(n110) );
  BUF_X1 U40 ( .A(n367), .Z(n111) );
  NAND2_X1 U41 ( .A1(n379), .A2(n386), .ZN(n445) );
  NOR2_X1 U42 ( .A1(opcode_i[14]), .A2(n376), .ZN(n367) );
  INV_X1 U43 ( .A(valid_i), .ZN(n286) );
  NOR2_X1 U44 ( .A1(n289), .A2(n391), .ZN(n374) );
  INV_X1 U45 ( .A(opcode_i[14]), .ZN(n386) );
  INV_X1 U46 ( .A(opcode_i[12]), .ZN(n164) );
  INV_X1 U47 ( .A(n380), .ZN(n447) );
  OAI21_X1 U48 ( .B1(n387), .B2(n386), .A(n380), .ZN(n442) );
  OAI21_X1 U49 ( .B1(n386), .B2(n371), .A(n370), .ZN(n365) );
  INV_X1 U50 ( .A(opcode_i[13]), .ZN(n147) );
  INV_X1 U51 ( .A(opcode_i[20]), .ZN(n211) );
  NOR2_X1 U52 ( .A1(n179), .A2(n96), .ZN(n109) );
  NOR2_X1 U53 ( .A1(n179), .A2(n97), .ZN(n108) );
  INV_X1 U54 ( .A(n188), .ZN(n107) );
  MUX2_X1 U55 ( .A(n107), .B(n108), .S(n311), .Z(n180) );
  MUX2_X1 U56 ( .A(n107), .B(n109), .S(n307), .Z(n177) );
  INV_X1 U57 ( .A(opcode_i[31]), .ZN(n113) );
  NAND3_X1 U58 ( .A1(csr_mcycle_q[2]), .A2(csr_mcycle_q[1]), .A3(
        csr_mcycle_q[0]), .ZN(n141) );
  NOR2_X1 U59 ( .A1(n86), .A2(n141), .ZN(n140) );
  NAND2_X1 U60 ( .A1(csr_mcycle_q[4]), .A2(n140), .ZN(n139) );
  NOR2_X1 U61 ( .A1(n95), .A2(n139), .ZN(n138) );
  NAND2_X1 U62 ( .A1(csr_mcycle_q[6]), .A2(n138), .ZN(n137) );
  NOR2_X1 U63 ( .A1(n94), .A2(n137), .ZN(n136) );
  NAND2_X1 U64 ( .A1(csr_mcycle_q[8]), .A2(n136), .ZN(n135) );
  NOR2_X1 U65 ( .A1(n93), .A2(n135), .ZN(n134) );
  NAND2_X1 U66 ( .A1(csr_mcycle_q[10]), .A2(n134), .ZN(n133) );
  NOR2_X1 U67 ( .A1(n92), .A2(n133), .ZN(n132) );
  NAND2_X1 U68 ( .A1(csr_mcycle_q[12]), .A2(n132), .ZN(n131) );
  NOR2_X1 U69 ( .A1(n91), .A2(n131), .ZN(n130) );
  NAND2_X1 U70 ( .A1(csr_mcycle_q[14]), .A2(n130), .ZN(n129) );
  NOR2_X1 U71 ( .A1(n90), .A2(n129), .ZN(n128) );
  NAND2_X1 U72 ( .A1(csr_mcycle_q[16]), .A2(n128), .ZN(n127) );
  NOR2_X1 U73 ( .A1(n89), .A2(n127), .ZN(n126) );
  NAND2_X1 U74 ( .A1(csr_mcycle_q[18]), .A2(n126), .ZN(n125) );
  NOR2_X1 U75 ( .A1(n88), .A2(n125), .ZN(n124) );
  NAND2_X1 U76 ( .A1(csr_mcycle_q[20]), .A2(n124), .ZN(n123) );
  NOR2_X1 U77 ( .A1(n87), .A2(n123), .ZN(n122) );
  NAND2_X1 U78 ( .A1(csr_mcycle_q[22]), .A2(n122), .ZN(n121) );
  NOR2_X1 U79 ( .A1(n102), .A2(n121), .ZN(n120) );
  NAND2_X1 U80 ( .A1(csr_mcycle_q[24]), .A2(n120), .ZN(n119) );
  NOR2_X1 U81 ( .A1(n101), .A2(n119), .ZN(n117) );
  NAND2_X1 U82 ( .A1(csr_mcycle_q[26]), .A2(n117), .ZN(n116) );
  NOR2_X1 U83 ( .A1(n100), .A2(n116), .ZN(n115) );
  NAND2_X1 U84 ( .A1(csr_mcycle_q[28]), .A2(n115), .ZN(n114) );
  NOR2_X1 U85 ( .A1(n99), .A2(n114), .ZN(n144) );
  XOR2_X1 U86 ( .A(csr_mcycle_q[30]), .B(n144), .Z(csr_mcycle_r[30]) );
  AOI21_X1 U87 ( .B1(n99), .B2(n114), .A(n144), .ZN(csr_mcycle_r[29]) );
  XOR2_X1 U88 ( .A(csr_mcycle_q[28]), .B(n115), .Z(csr_mcycle_r[28]) );
  AOI21_X1 U89 ( .B1(n100), .B2(n116), .A(n115), .ZN(csr_mcycle_r[27]) );
  XOR2_X1 U90 ( .A(csr_mcycle_q[26]), .B(n117), .Z(csr_mcycle_r[26]) );
  AOI21_X1 U91 ( .B1(n101), .B2(n119), .A(n117), .ZN(csr_mcycle_r[25]) );
  XOR2_X1 U92 ( .A(csr_mcycle_q[24]), .B(n120), .Z(csr_mcycle_r[24]) );
  AOI21_X1 U93 ( .B1(n102), .B2(n121), .A(n120), .ZN(csr_mcycle_r[23]) );
  XOR2_X1 U94 ( .A(csr_mcycle_q[22]), .B(n122), .Z(csr_mcycle_r[22]) );
  AOI21_X1 U95 ( .B1(n87), .B2(n123), .A(n122), .ZN(csr_mcycle_r[21]) );
  XOR2_X1 U96 ( .A(csr_mcycle_q[20]), .B(n124), .Z(csr_mcycle_r[20]) );
  AOI21_X1 U97 ( .B1(n88), .B2(n125), .A(n124), .ZN(csr_mcycle_r[19]) );
  XOR2_X1 U98 ( .A(csr_mcycle_q[18]), .B(n126), .Z(csr_mcycle_r[18]) );
  AOI21_X1 U99 ( .B1(n89), .B2(n127), .A(n126), .ZN(csr_mcycle_r[17]) );
  XOR2_X1 U100 ( .A(csr_mcycle_q[16]), .B(n128), .Z(csr_mcycle_r[16]) );
  AOI21_X1 U101 ( .B1(n90), .B2(n129), .A(n128), .ZN(csr_mcycle_r[15]) );
  XOR2_X1 U102 ( .A(csr_mcycle_q[14]), .B(n130), .Z(csr_mcycle_r[14]) );
  AOI21_X1 U103 ( .B1(n91), .B2(n131), .A(n130), .ZN(csr_mcycle_r[13]) );
  XOR2_X1 U104 ( .A(csr_mcycle_q[12]), .B(n132), .Z(csr_mcycle_r[12]) );
  AOI21_X1 U105 ( .B1(n92), .B2(n133), .A(n132), .ZN(csr_mcycle_r[11]) );
  XOR2_X1 U106 ( .A(csr_mcycle_q[10]), .B(n134), .Z(csr_mcycle_r[10]) );
  AOI21_X1 U107 ( .B1(n93), .B2(n135), .A(n134), .ZN(csr_mcycle_r[9]) );
  XOR2_X1 U108 ( .A(csr_mcycle_q[8]), .B(n136), .Z(csr_mcycle_r[8]) );
  AOI21_X1 U109 ( .B1(n94), .B2(n137), .A(n136), .ZN(csr_mcycle_r[7]) );
  XOR2_X1 U110 ( .A(csr_mcycle_q[6]), .B(n138), .Z(csr_mcycle_r[6]) );
  AOI21_X1 U111 ( .B1(n95), .B2(n139), .A(n138), .ZN(csr_mcycle_r[5]) );
  XOR2_X1 U112 ( .A(csr_mcycle_q[4]), .B(n140), .Z(csr_mcycle_r[4]) );
  NOR2_X1 U113 ( .A1(n98), .A2(n85), .ZN(n143) );
  OAI21_X1 U114 ( .B1(csr_mcycle_q[2]), .B2(n143), .A(n141), .ZN(n142) );
  NAND2_X1 U115 ( .A1(csr_mcycle_q[30]), .A2(n144), .ZN(n145) );
  XNOR2_X1 U116 ( .A(csr_mcycle_q[31]), .B(n145), .ZN(csr_mcycle_r[31]) );
  NOR2_X1 U117 ( .A1(opcode_i[3]), .A2(opcode_i[2]), .ZN(n171) );
  NAND4_X1 U118 ( .A1(opcode_i[5]), .A2(opcode_i[4]), .A3(opcode_i[6]), .A4(
        n171), .ZN(n153) );
  OR2_X1 U119 ( .A1(exception_o), .A2(n153), .ZN(n163) );
  NOR3_X1 U120 ( .A1(n147), .A2(n164), .A3(n163), .ZN(n290) );
  INV_X1 U121 ( .A(n290), .ZN(n179) );
  NOR2_X1 U122 ( .A1(n179), .A2(n103), .ZN(n156) );
  AOI22_X1 U123 ( .A1(opcode_i[14]), .A2(opcode_i[15]), .B1(rs1_val_i[0]), 
        .B2(n386), .ZN(n299) );
  AOI221_X1 U124 ( .B1(opcode_i[13]), .B2(opcode_i[12]), .C1(n147), .C2(n164), 
        .A(n163), .ZN(n288) );
  INV_X1 U125 ( .A(opcode_i[30]), .ZN(n201) );
  NAND2_X1 U126 ( .A1(n211), .A2(n201), .ZN(n157) );
  INV_X1 U127 ( .A(opcode_i[21]), .ZN(n148) );
  NOR3_X1 U128 ( .A1(opcode_i[25]), .A2(opcode_i[24]), .A3(opcode_i[23]), .ZN(
        n191) );
  NAND2_X1 U129 ( .A1(n191), .A2(opcode_i[28]), .ZN(n159) );
  NAND2_X1 U130 ( .A1(valid_i), .A2(opcode_i[29]), .ZN(n197) );
  NOR3_X1 U131 ( .A1(opcode_i[31]), .A2(n159), .A3(n197), .ZN(n208) );
  NAND2_X1 U132 ( .A1(n288), .A2(n256), .ZN(n188) );
  INV_X1 U133 ( .A(n299), .ZN(n296) );
  NOR2_X1 U134 ( .A1(opcode_i[26]), .A2(opcode_i[27]), .ZN(n193) );
  NOR2_X1 U135 ( .A1(opcode_i[21]), .A2(opcode_i[22]), .ZN(n200) );
  NAND2_X1 U136 ( .A1(n193), .A2(n200), .ZN(n189) );
  NOR2_X1 U137 ( .A1(opcode_i[30]), .A2(n189), .ZN(n209) );
  OR4_X1 U138 ( .A1(opcode_i[10]), .A2(opcode_i[11]), .A3(opcode_i[14]), .A4(
        opcode_i[12]), .ZN(n152) );
  NOR4_X1 U139 ( .A1(opcode_i[13]), .A2(opcode_i[17]), .A3(opcode_i[16]), .A4(
        opcode_i[18]), .ZN(n150) );
  NOR4_X1 U140 ( .A1(opcode_i[7]), .A2(opcode_i[19]), .A3(opcode_i[8]), .A4(
        opcode_i[9]), .ZN(n149) );
  NAND2_X1 U141 ( .A1(n150), .A2(n149), .ZN(n151) );
  NOR4_X1 U142 ( .A1(opcode_i[15]), .A2(n153), .A3(n152), .A4(n151), .ZN(n162)
         );
  INV_X1 U143 ( .A(n162), .ZN(n154) );
  NOR4_X1 U144 ( .A1(opcode_i[31]), .A2(opcode_i[29]), .A3(opcode_i[28]), .A4(
        n154), .ZN(n155) );
  NAND3_X1 U145 ( .A1(n191), .A2(n209), .A3(n155), .ZN(n165) );
  NOR3_X1 U146 ( .A1(excpn_invalid_inst_i), .A2(n286), .A3(n165), .ZN(n181) );
  AOI221_X1 U147 ( .B1(n156), .B2(n299), .C1(n107), .C2(n296), .A(n181), .ZN(
        n167) );
  INV_X1 U148 ( .A(n157), .ZN(n158) );
  NAND2_X1 U149 ( .A1(opcode_i[29]), .A2(n158), .ZN(n160) );
  NOR4_X1 U150 ( .A1(opcode_i[31]), .A2(opcode_i[22]), .A3(n160), .A4(n159), 
        .ZN(n161) );
  NAND4_X1 U151 ( .A1(n162), .A2(opcode_i[21]), .A3(n193), .A4(n161), .ZN(n278) );
  NOR2_X1 U152 ( .A1(n164), .A2(n163), .ZN(n293) );
  NAND3_X1 U153 ( .A1(n278), .A2(n256), .A3(n293), .ZN(n166) );
  INV_X1 U154 ( .A(n165), .ZN(n169) );
  NOR2_X1 U155 ( .A1(exception_o), .A2(n169), .ZN(n289) );
  NAND2_X1 U156 ( .A1(n166), .A2(n289), .ZN(n168) );
  NAND2_X1 U157 ( .A1(valid_i), .A2(n168), .ZN(n185) );
  NAND2_X1 U158 ( .A1(n118), .A2(n185), .ZN(n182) );
  OAI22_X1 U159 ( .A1(rst_i), .A2(n167), .B1(n182), .B2(n103), .ZN(N818) );
  AOI22_X1 U160 ( .A1(opcode_i[14]), .A2(opcode_i[16]), .B1(rs1_val_i[1]), 
        .B2(n386), .ZN(n303) );
  INV_X1 U161 ( .A(n303), .ZN(n300) );
  OAI21_X1 U162 ( .B1(n179), .B2(n300), .A(n168), .ZN(n174) );
  OR2_X1 U163 ( .A1(excpn_invalid_inst_i), .A2(n169), .ZN(n176) );
  INV_X1 U164 ( .A(opcode_i[4]), .ZN(n170) );
  NAND4_X1 U165 ( .A1(opcode_i[5]), .A2(n171), .A3(excpn_lsu_align_i), .A4(
        n170), .ZN(n172) );
  OAI22_X1 U166 ( .A1(n303), .A2(n188), .B1(opcode_i[6]), .B2(n172), .ZN(n173)
         );
  AOI211_X1 U167 ( .C1(csr_mcause_q[1]), .C2(n174), .A(n176), .B(n173), .ZN(
        n175) );
  AOI221_X1 U168 ( .B1(valid_i), .B2(n175), .C1(n286), .C2(n105), .A(rst_i), 
        .ZN(N819) );
  NOR2_X1 U169 ( .A1(n289), .A2(n176), .ZN(n184) );
  AOI22_X1 U171 ( .A1(opcode_i[14]), .A2(opcode_i[17]), .B1(rs1_val_i[2]), 
        .B2(n386), .ZN(n307) );
  INV_X1 U172 ( .A(n307), .ZN(n304) );
  AOI21_X1 U173 ( .B1(excpn_lsu_align_i), .B2(n184), .A(n177), .ZN(n178) );
  OAI22_X1 U174 ( .A1(rst_i), .A2(n178), .B1(n96), .B2(n182), .ZN(N820) );
  AOI22_X1 U175 ( .A1(opcode_i[14]), .A2(opcode_i[18]), .B1(rs1_val_i[3]), 
        .B2(n386), .ZN(n311) );
  INV_X1 U176 ( .A(n311), .ZN(n308) );
  AOI21_X1 U177 ( .B1(n181), .B2(n211), .A(n180), .ZN(n183) );
  OAI22_X1 U178 ( .A1(rst_i), .A2(n183), .B1(n97), .B2(n182), .ZN(N821) );
  NAND2_X1 U179 ( .A1(rs1_val_i[31]), .A2(n386), .ZN(n449) );
  INV_X1 U180 ( .A(n184), .ZN(n187) );
  AOI21_X1 U181 ( .B1(n290), .B2(n449), .A(n185), .ZN(n186) );
  OAI222_X1 U182 ( .A1(n188), .A2(n449), .B1(n187), .B2(excpn_lsu_align_i), 
        .C1(n104), .C2(n186), .ZN(csr_mcause_r_31_) );
  NOR4_X1 U183 ( .A1(opcode_i[29]), .A2(opcode_i[28]), .A3(n201), .A4(n189), 
        .ZN(n190) );
  NAND4_X1 U184 ( .A1(valid_i), .A2(opcode_i[31]), .A3(n191), .A4(n190), .ZN(
        n259) );
  INV_X1 U185 ( .A(opcode_i[25]), .ZN(n192) );
  NAND3_X1 U186 ( .A1(n193), .A2(opcode_i[24]), .A3(n192), .ZN(n196) );
  NOR3_X1 U187 ( .A1(opcode_i[20]), .A2(opcode_i[23]), .A3(n113), .ZN(n194) );
  NAND4_X1 U188 ( .A1(opcode_i[30]), .A2(opcode_i[28]), .A3(opcode_i[22]), 
        .A4(n194), .ZN(n195) );
  NOR4_X1 U189 ( .A1(opcode_i[21]), .A2(n197), .A3(n196), .A4(n195), .ZN(n273)
         );
  AOI22_X1 U190 ( .A1(n256), .A2(csr_mcause_q[0]), .B1(n82), .B2(cpu_id_i[0]), 
        .ZN(n203) );
  INV_X1 U191 ( .A(n198), .ZN(n199) );
  NAND4_X1 U192 ( .A1(n201), .A2(opcode_i[20]), .A3(n200), .A4(n199), .ZN(n271) );
  AOI22_X1 U193 ( .A1(n292), .A2(csr_mepc_o[0]), .B1(n276), .B2(csr_sr_q[0]), 
        .ZN(n202) );
  OAI211_X1 U194 ( .C1(n85), .C2(n259), .A(n203), .B(n202), .ZN(csr_rdata_o[0]) );
  AOI22_X1 U195 ( .A1(csr_mcycle_q[10]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[10]), .ZN(n205) );
  AOI22_X1 U196 ( .A1(n276), .A2(csr_sr_q[10]), .B1(n82), .B2(cpu_id_i[10]), 
        .ZN(n204) );
  NAND2_X1 U197 ( .A1(n205), .A2(n204), .ZN(csr_rdata_o[10]) );
  AOI22_X1 U198 ( .A1(csr_mcycle_q[11]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[11]), .ZN(n207) );
  AOI22_X1 U199 ( .A1(n276), .A2(csr_sr_q[11]), .B1(n82), .B2(cpu_id_i[11]), 
        .ZN(n206) );
  NAND2_X1 U200 ( .A1(n207), .A2(n206), .ZN(csr_rdata_o[11]) );
  NAND2_X1 U201 ( .A1(n209), .A2(n208), .ZN(n210) );
  NOR2_X1 U202 ( .A1(n211), .A2(n210), .ZN(n268) );
  AOI21_X1 U203 ( .B1(n82), .B2(cpu_id_i[12]), .A(n268), .ZN(n213) );
  AOI22_X1 U204 ( .A1(csr_mcycle_q[12]), .A2(n272), .B1(n276), .B2(
        csr_sr_q[12]), .ZN(n212) );
  OAI211_X1 U205 ( .C1(n64), .C2(n271), .A(n213), .B(n212), .ZN(
        csr_rdata_o[12]) );
  AOI22_X1 U206 ( .A1(csr_mcycle_q[13]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[13]), .ZN(n215) );
  AOI22_X1 U207 ( .A1(n276), .A2(csr_sr_q[13]), .B1(n82), .B2(cpu_id_i[13]), 
        .ZN(n214) );
  NAND2_X1 U208 ( .A1(n215), .A2(n214), .ZN(csr_rdata_o[13]) );
  AOI22_X1 U209 ( .A1(csr_mcycle_q[14]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[14]), .ZN(n217) );
  AOI22_X1 U210 ( .A1(n276), .A2(csr_sr_q[14]), .B1(n82), .B2(cpu_id_i[14]), 
        .ZN(n216) );
  NAND2_X1 U211 ( .A1(n217), .A2(n216), .ZN(csr_rdata_o[14]) );
  AOI22_X1 U212 ( .A1(csr_mcycle_q[15]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[15]), .ZN(n219) );
  AOI22_X1 U213 ( .A1(n276), .A2(csr_sr_q[15]), .B1(n82), .B2(cpu_id_i[15]), 
        .ZN(n218) );
  NAND2_X1 U214 ( .A1(n219), .A2(n218), .ZN(csr_rdata_o[15]) );
  AOI22_X1 U215 ( .A1(csr_mcycle_q[16]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[16]), .ZN(n221) );
  AOI22_X1 U216 ( .A1(n276), .A2(csr_sr_q[16]), .B1(n82), .B2(cpu_id_i[16]), 
        .ZN(n220) );
  NAND2_X1 U217 ( .A1(n221), .A2(n220), .ZN(csr_rdata_o[16]) );
  AOI22_X1 U218 ( .A1(csr_mcycle_q[17]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[17]), .ZN(n223) );
  AOI22_X1 U219 ( .A1(n276), .A2(csr_sr_q[17]), .B1(n82), .B2(cpu_id_i[17]), 
        .ZN(n222) );
  NAND2_X1 U220 ( .A1(n223), .A2(n222), .ZN(csr_rdata_o[17]) );
  AOI22_X1 U221 ( .A1(csr_mcycle_q[18]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[18]), .ZN(n225) );
  AOI22_X1 U222 ( .A1(n276), .A2(csr_sr_q[18]), .B1(n82), .B2(cpu_id_i[18]), 
        .ZN(n224) );
  NAND2_X1 U223 ( .A1(n225), .A2(n224), .ZN(csr_rdata_o[18]) );
  AOI22_X1 U224 ( .A1(csr_mcycle_q[19]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[19]), .ZN(n227) );
  AOI22_X1 U225 ( .A1(n276), .A2(csr_sr_q[19]), .B1(n82), .B2(cpu_id_i[19]), 
        .ZN(n226) );
  NAND2_X1 U226 ( .A1(n227), .A2(n226), .ZN(csr_rdata_o[19]) );
  AOI22_X1 U227 ( .A1(csr_mcause_q[1]), .A2(n256), .B1(n82), .B2(cpu_id_i[1]), 
        .ZN(n229) );
  AOI22_X1 U228 ( .A1(csr_mcycle_q[1]), .A2(n272), .B1(n276), .B2(csr_sr_q[1]), 
        .ZN(n228) );
  OAI211_X1 U229 ( .C1(n75), .C2(n271), .A(n229), .B(n228), .ZN(csr_rdata_o[1]) );
  AOI22_X1 U230 ( .A1(csr_mcycle_q[20]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[20]), .ZN(n231) );
  AOI22_X1 U231 ( .A1(n276), .A2(csr_sr_q[20]), .B1(n82), .B2(cpu_id_i[20]), 
        .ZN(n230) );
  NAND2_X1 U232 ( .A1(n231), .A2(n230), .ZN(csr_rdata_o[20]) );
  AOI22_X1 U233 ( .A1(csr_mcycle_q[21]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[21]), .ZN(n233) );
  AOI22_X1 U234 ( .A1(n276), .A2(csr_sr_q[21]), .B1(n82), .B2(cpu_id_i[21]), 
        .ZN(n232) );
  NAND2_X1 U235 ( .A1(n233), .A2(n232), .ZN(csr_rdata_o[21]) );
  AOI22_X1 U236 ( .A1(csr_mcycle_q[22]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[22]), .ZN(n235) );
  AOI22_X1 U237 ( .A1(n276), .A2(csr_sr_q[22]), .B1(n82), .B2(cpu_id_i[22]), 
        .ZN(n234) );
  NAND2_X1 U238 ( .A1(n235), .A2(n234), .ZN(csr_rdata_o[22]) );
  AOI22_X1 U239 ( .A1(csr_mcycle_q[23]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[23]), .ZN(n237) );
  AOI22_X1 U240 ( .A1(n276), .A2(csr_sr_q[23]), .B1(n82), .B2(cpu_id_i[23]), 
        .ZN(n236) );
  NAND2_X1 U241 ( .A1(n237), .A2(n236), .ZN(csr_rdata_o[23]) );
  AOI22_X1 U242 ( .A1(csr_mcycle_q[24]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[24]), .ZN(n239) );
  AOI22_X1 U243 ( .A1(n276), .A2(csr_sr_q[24]), .B1(n82), .B2(cpu_id_i[24]), 
        .ZN(n238) );
  NAND2_X1 U244 ( .A1(n239), .A2(n238), .ZN(csr_rdata_o[24]) );
  AOI22_X1 U245 ( .A1(csr_mcycle_q[25]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[25]), .ZN(n241) );
  AOI22_X1 U246 ( .A1(n276), .A2(csr_sr_q[25]), .B1(n82), .B2(cpu_id_i[25]), 
        .ZN(n240) );
  NAND2_X1 U247 ( .A1(n241), .A2(n240), .ZN(csr_rdata_o[25]) );
  AOI22_X1 U248 ( .A1(csr_mcycle_q[26]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[26]), .ZN(n243) );
  AOI22_X1 U249 ( .A1(n276), .A2(csr_sr_q[26]), .B1(n82), .B2(cpu_id_i[26]), 
        .ZN(n242) );
  NAND2_X1 U250 ( .A1(n243), .A2(n242), .ZN(csr_rdata_o[26]) );
  AOI22_X1 U251 ( .A1(csr_mcycle_q[27]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[27]), .ZN(n245) );
  AOI22_X1 U252 ( .A1(n276), .A2(csr_sr_q[27]), .B1(n82), .B2(cpu_id_i[27]), 
        .ZN(n244) );
  NAND2_X1 U253 ( .A1(n245), .A2(n244), .ZN(csr_rdata_o[27]) );
  AOI22_X1 U254 ( .A1(csr_mcycle_q[28]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[28]), .ZN(n247) );
  AOI22_X1 U255 ( .A1(n276), .A2(csr_sr_q[28]), .B1(n82), .B2(cpu_id_i[28]), 
        .ZN(n246) );
  NAND2_X1 U256 ( .A1(n247), .A2(n246), .ZN(csr_rdata_o[28]) );
  AOI22_X1 U257 ( .A1(csr_mcycle_q[29]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[29]), .ZN(n249) );
  AOI22_X1 U258 ( .A1(n276), .A2(csr_sr_q[29]), .B1(n82), .B2(cpu_id_i[29]), 
        .ZN(n248) );
  NAND2_X1 U259 ( .A1(n249), .A2(n248), .ZN(csr_rdata_o[29]) );
  AOI22_X1 U260 ( .A1(n256), .A2(csr_mcause_q[2]), .B1(n82), .B2(cpu_id_i[2]), 
        .ZN(n251) );
  AOI22_X1 U261 ( .A1(csr_mcycle_q[2]), .A2(n272), .B1(n276), .B2(csr_sr_q[2]), 
        .ZN(n250) );
  OAI211_X1 U262 ( .C1(n74), .C2(n271), .A(n251), .B(n250), .ZN(csr_rdata_o[2]) );
  AOI21_X1 U263 ( .B1(n82), .B2(cpu_id_i[30]), .A(n268), .ZN(n253) );
  AOI22_X1 U264 ( .A1(csr_mcycle_q[30]), .A2(n272), .B1(n276), .B2(
        csr_sr_q[30]), .ZN(n252) );
  OAI211_X1 U265 ( .C1(n46), .C2(n271), .A(n253), .B(n252), .ZN(
        csr_rdata_o[30]) );
  AOI22_X1 U266 ( .A1(n256), .A2(csr_mcause_q[31]), .B1(n82), .B2(cpu_id_i[31]), .ZN(n255) );
  AOI22_X1 U267 ( .A1(csr_mcycle_q[31]), .A2(n272), .B1(n276), .B2(
        csr_sr_q[31]), .ZN(n254) );
  OAI211_X1 U268 ( .C1(n45), .C2(n271), .A(n255), .B(n254), .ZN(
        csr_rdata_o[31]) );
  AOI22_X1 U269 ( .A1(n256), .A2(csr_mcause_q[3]), .B1(n82), .B2(cpu_id_i[3]), 
        .ZN(n258) );
  AOI22_X1 U270 ( .A1(csr_sr_q[3]), .A2(n276), .B1(n292), .B2(csr_mepc_o[3]), 
        .ZN(n257) );
  OAI211_X1 U271 ( .C1(n86), .C2(n259), .A(n258), .B(n257), .ZN(csr_rdata_o[3]) );
  AOI22_X1 U272 ( .A1(csr_mcycle_q[4]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[4]), .ZN(n261) );
  AOI22_X1 U273 ( .A1(n276), .A2(csr_sr_q[4]), .B1(n82), .B2(cpu_id_i[4]), 
        .ZN(n260) );
  NAND2_X1 U274 ( .A1(n261), .A2(n260), .ZN(csr_rdata_o[4]) );
  AOI22_X1 U275 ( .A1(csr_mcycle_q[5]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[5]), .ZN(n263) );
  AOI22_X1 U276 ( .A1(n276), .A2(csr_sr_q[5]), .B1(n82), .B2(cpu_id_i[5]), 
        .ZN(n262) );
  NAND2_X1 U277 ( .A1(n263), .A2(n262), .ZN(csr_rdata_o[5]) );
  AOI22_X1 U278 ( .A1(csr_mcycle_q[6]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[6]), .ZN(n265) );
  AOI22_X1 U279 ( .A1(n276), .A2(csr_sr_q[6]), .B1(n82), .B2(cpu_id_i[6]), 
        .ZN(n264) );
  NAND2_X1 U280 ( .A1(n265), .A2(n264), .ZN(csr_rdata_o[6]) );
  AOI22_X1 U281 ( .A1(csr_mcycle_q[7]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[7]), .ZN(n267) );
  AOI22_X1 U282 ( .A1(n276), .A2(csr_sr_q[7]), .B1(n82), .B2(cpu_id_i[7]), 
        .ZN(n266) );
  NAND2_X1 U283 ( .A1(n267), .A2(n266), .ZN(csr_rdata_o[7]) );
  AOI22_X1 U284 ( .A1(csr_mcycle_q[8]), .A2(n272), .B1(n82), .B2(cpu_id_i[8]), 
        .ZN(n270) );
  AOI21_X1 U285 ( .B1(csr_sr_q[8]), .B2(n276), .A(n268), .ZN(n269) );
  OAI211_X1 U286 ( .C1(n68), .C2(n271), .A(n270), .B(n269), .ZN(csr_rdata_o[8]) );
  AOI22_X1 U287 ( .A1(csr_mcycle_q[9]), .A2(n272), .B1(n292), .B2(
        csr_mepc_o[9]), .ZN(n275) );
  AOI22_X1 U288 ( .A1(n276), .A2(csr_sr_q[9]), .B1(n82), .B2(cpu_id_i[9]), 
        .ZN(n274) );
  NAND2_X1 U289 ( .A1(n275), .A2(n274), .ZN(csr_rdata_o[9]) );
  NAND3_X1 U290 ( .A1(n118), .A2(n288), .A3(n276), .ZN(n450) );
  NAND2_X1 U291 ( .A1(n293), .A2(n276), .ZN(n279) );
  NAND2_X1 U292 ( .A1(n118), .A2(n279), .ZN(n380) );
  NAND2_X1 U293 ( .A1(n118), .A2(n290), .ZN(n387) );
  OAI221_X1 U294 ( .B1(n447), .B2(n299), .C1(n447), .C2(n446), .A(csr_sr_q[0]), 
        .ZN(n277) );
  OAI21_X1 U295 ( .B1(n299), .B2(n450), .A(n277), .ZN(n623) );
  NOR2_X1 U296 ( .A1(n286), .A2(rst_i), .ZN(n401) );
  INV_X1 U297 ( .A(n289), .ZN(n389) );
  NOR2_X1 U298 ( .A1(n278), .A2(n389), .ZN(n388) );
  NAND3_X1 U299 ( .A1(n401), .A2(csr_sr_q[7]), .A3(n388), .ZN(n283) );
  NAND2_X1 U300 ( .A1(n289), .A2(n278), .ZN(n400) );
  INV_X1 U301 ( .A(n400), .ZN(n280) );
  OAI221_X1 U302 ( .B1(n286), .B2(n280), .C1(n286), .C2(n279), .A(n118), .ZN(
        n385) );
  OAI21_X1 U303 ( .B1(n387), .B2(n308), .A(n385), .ZN(n281) );
  INV_X1 U304 ( .A(n450), .ZN(n379) );
  AOI22_X1 U305 ( .A1(csr_sr_q[3]), .A2(n281), .B1(n379), .B2(n308), .ZN(n282)
         );
  NAND2_X1 U306 ( .A1(n283), .A2(n282), .ZN(n622) );
  OAI221_X1 U307 ( .B1(n447), .B2(n307), .C1(n447), .C2(n446), .A(csr_sr_q[2]), 
        .ZN(n284) );
  OAI21_X1 U308 ( .B1(n307), .B2(n450), .A(n284), .ZN(n621) );
  OAI221_X1 U309 ( .B1(n447), .B2(n303), .C1(n447), .C2(n446), .A(csr_sr_q[1]), 
        .ZN(n285) );
  OAI21_X1 U310 ( .B1(n303), .B2(n450), .A(n285), .ZN(n620) );
  OAI21_X1 U311 ( .B1(n388), .B2(n286), .A(n118), .ZN(n287) );
  INV_X1 U312 ( .A(n287), .ZN(n294) );
  NOR2_X1 U313 ( .A1(rst_i), .A2(n294), .ZN(n291) );
  NAND3_X1 U314 ( .A1(n291), .A2(n292), .A3(n288), .ZN(n376) );
  INV_X1 U315 ( .A(n401), .ZN(n391) );
  NAND2_X1 U316 ( .A1(n291), .A2(n290), .ZN(n371) );
  AOI21_X1 U317 ( .B1(n293), .B2(n292), .A(n400), .ZN(n295) );
  AOI21_X1 U318 ( .B1(n295), .B2(n118), .A(n294), .ZN(n370) );
  OAI21_X1 U319 ( .B1(n371), .B2(n296), .A(n370), .ZN(n297) );
  AOI22_X1 U320 ( .A1(n374), .A2(pc_i[0]), .B1(csr_mepc_o[0]), .B2(n297), .ZN(
        n298) );
  OAI21_X1 U321 ( .B1(n299), .B2(n376), .A(n298), .ZN(n619) );
  OAI21_X1 U322 ( .B1(n371), .B2(n300), .A(n370), .ZN(n301) );
  AOI22_X1 U323 ( .A1(n374), .A2(pc_i[1]), .B1(csr_mepc_o[1]), .B2(n301), .ZN(
        n302) );
  OAI21_X1 U324 ( .B1(n303), .B2(n376), .A(n302), .ZN(n618) );
  OAI21_X1 U325 ( .B1(n371), .B2(n304), .A(n370), .ZN(n305) );
  AOI22_X1 U326 ( .A1(n374), .A2(pc_i[2]), .B1(csr_mepc_o[2]), .B2(n305), .ZN(
        n306) );
  OAI21_X1 U327 ( .B1(n307), .B2(n376), .A(n306), .ZN(n617) );
  OAI21_X1 U328 ( .B1(n371), .B2(n308), .A(n370), .ZN(n309) );
  AOI22_X1 U329 ( .A1(n112), .A2(pc_i[3]), .B1(csr_mepc_o[3]), .B2(n309), .ZN(
        n310) );
  OAI21_X1 U330 ( .B1(n311), .B2(n376), .A(n310), .ZN(n616) );
  AOI22_X1 U331 ( .A1(opcode_i[14]), .A2(opcode_i[19]), .B1(rs1_val_i[4]), 
        .B2(n386), .ZN(n378) );
  INV_X1 U332 ( .A(n378), .ZN(n312) );
  OAI21_X1 U333 ( .B1(n371), .B2(n312), .A(n370), .ZN(n313) );
  AOI22_X1 U334 ( .A1(n112), .A2(pc_i[4]), .B1(csr_mepc_o[4]), .B2(n313), .ZN(
        n314) );
  OAI21_X1 U335 ( .B1(n378), .B2(n376), .A(n314), .ZN(n615) );
  INV_X1 U336 ( .A(rs1_val_i[5]), .ZN(n382) );
  AOI21_X1 U337 ( .B1(n366), .B2(n382), .A(n110), .ZN(n316) );
  AOI22_X1 U338 ( .A1(rs1_val_i[5]), .A2(n367), .B1(n374), .B2(pc_i[5]), .ZN(
        n315) );
  OAI21_X1 U339 ( .B1(n71), .B2(n316), .A(n315), .ZN(n614) );
  INV_X1 U340 ( .A(rs1_val_i[6]), .ZN(n384) );
  AOI21_X1 U341 ( .B1(n366), .B2(n384), .A(n110), .ZN(n318) );
  AOI22_X1 U342 ( .A1(n111), .A2(rs1_val_i[6]), .B1(n112), .B2(pc_i[6]), .ZN(
        n317) );
  OAI21_X1 U343 ( .B1(n70), .B2(n318), .A(n317), .ZN(n613) );
  INV_X1 U344 ( .A(rs1_val_i[7]), .ZN(n393) );
  AOI21_X1 U345 ( .B1(n366), .B2(n393), .A(n110), .ZN(n320) );
  AOI22_X1 U346 ( .A1(n367), .A2(rs1_val_i[7]), .B1(n112), .B2(pc_i[7]), .ZN(
        n319) );
  OAI21_X1 U347 ( .B1(n69), .B2(n320), .A(n319), .ZN(n612) );
  INV_X1 U348 ( .A(rs1_val_i[8]), .ZN(n395) );
  AOI21_X1 U349 ( .B1(n366), .B2(n395), .A(n110), .ZN(n322) );
  AOI22_X1 U350 ( .A1(n367), .A2(rs1_val_i[8]), .B1(n112), .B2(pc_i[8]), .ZN(
        n321) );
  OAI21_X1 U351 ( .B1(n68), .B2(n322), .A(n321), .ZN(n611) );
  INV_X1 U352 ( .A(rs1_val_i[9]), .ZN(n397) );
  AOI21_X1 U353 ( .B1(n366), .B2(n397), .A(n110), .ZN(n324) );
  AOI22_X1 U354 ( .A1(n367), .A2(rs1_val_i[9]), .B1(n374), .B2(pc_i[9]), .ZN(
        n323) );
  OAI21_X1 U355 ( .B1(n67), .B2(n324), .A(n323), .ZN(n610) );
  INV_X1 U356 ( .A(rs1_val_i[10]), .ZN(n399) );
  AOI21_X1 U357 ( .B1(n366), .B2(n399), .A(n110), .ZN(n326) );
  AOI22_X1 U358 ( .A1(n367), .A2(rs1_val_i[10]), .B1(n112), .B2(pc_i[10]), 
        .ZN(n325) );
  OAI21_X1 U359 ( .B1(n66), .B2(n326), .A(n325), .ZN(n609) );
  INV_X1 U360 ( .A(rs1_val_i[11]), .ZN(n403) );
  AOI21_X1 U361 ( .B1(n366), .B2(n403), .A(n110), .ZN(n328) );
  AOI22_X1 U362 ( .A1(n367), .A2(rs1_val_i[11]), .B1(n374), .B2(pc_i[11]), 
        .ZN(n327) );
  OAI21_X1 U363 ( .B1(n65), .B2(n328), .A(n327), .ZN(n608) );
  INV_X1 U364 ( .A(rs1_val_i[12]), .ZN(n407) );
  AOI21_X1 U365 ( .B1(n366), .B2(n407), .A(n110), .ZN(n330) );
  AOI22_X1 U366 ( .A1(n367), .A2(rs1_val_i[12]), .B1(n374), .B2(pc_i[12]), 
        .ZN(n329) );
  OAI21_X1 U367 ( .B1(n64), .B2(n330), .A(n329), .ZN(n607) );
  INV_X1 U368 ( .A(rs1_val_i[13]), .ZN(n409) );
  AOI21_X1 U369 ( .B1(n366), .B2(n409), .A(n110), .ZN(n332) );
  AOI22_X1 U370 ( .A1(n111), .A2(rs1_val_i[13]), .B1(n112), .B2(pc_i[13]), 
        .ZN(n331) );
  OAI21_X1 U371 ( .B1(n63), .B2(n332), .A(n331), .ZN(n606) );
  INV_X1 U372 ( .A(rs1_val_i[14]), .ZN(n411) );
  AOI21_X1 U373 ( .B1(n366), .B2(n411), .A(n110), .ZN(n334) );
  AOI22_X1 U374 ( .A1(n367), .A2(rs1_val_i[14]), .B1(n112), .B2(pc_i[14]), 
        .ZN(n333) );
  OAI21_X1 U375 ( .B1(n62), .B2(n334), .A(n333), .ZN(n605) );
  INV_X1 U376 ( .A(rs1_val_i[15]), .ZN(n413) );
  AOI21_X1 U377 ( .B1(n366), .B2(n413), .A(n110), .ZN(n336) );
  AOI22_X1 U378 ( .A1(n367), .A2(rs1_val_i[15]), .B1(n112), .B2(pc_i[15]), 
        .ZN(n335) );
  OAI21_X1 U379 ( .B1(n61), .B2(n336), .A(n335), .ZN(n604) );
  INV_X1 U380 ( .A(rs1_val_i[16]), .ZN(n415) );
  AOI21_X1 U381 ( .B1(n366), .B2(n415), .A(n110), .ZN(n338) );
  AOI22_X1 U382 ( .A1(n367), .A2(rs1_val_i[16]), .B1(n112), .B2(pc_i[16]), 
        .ZN(n337) );
  OAI21_X1 U383 ( .B1(n60), .B2(n338), .A(n337), .ZN(n603) );
  INV_X1 U384 ( .A(rs1_val_i[17]), .ZN(n417) );
  AOI21_X1 U385 ( .B1(n366), .B2(n417), .A(n365), .ZN(n340) );
  AOI22_X1 U386 ( .A1(n367), .A2(rs1_val_i[17]), .B1(n112), .B2(pc_i[17]), 
        .ZN(n339) );
  OAI21_X1 U387 ( .B1(n59), .B2(n340), .A(n339), .ZN(n602) );
  INV_X1 U388 ( .A(rs1_val_i[18]), .ZN(n419) );
  AOI21_X1 U389 ( .B1(n366), .B2(n419), .A(n365), .ZN(n342) );
  AOI22_X1 U390 ( .A1(n367), .A2(rs1_val_i[18]), .B1(n112), .B2(pc_i[18]), 
        .ZN(n341) );
  OAI21_X1 U391 ( .B1(n58), .B2(n342), .A(n341), .ZN(n601) );
  INV_X1 U392 ( .A(rs1_val_i[19]), .ZN(n421) );
  AOI21_X1 U393 ( .B1(n366), .B2(n421), .A(n365), .ZN(n344) );
  AOI22_X1 U394 ( .A1(n111), .A2(rs1_val_i[19]), .B1(n112), .B2(pc_i[19]), 
        .ZN(n343) );
  OAI21_X1 U395 ( .B1(n57), .B2(n344), .A(n343), .ZN(n600) );
  INV_X1 U396 ( .A(rs1_val_i[20]), .ZN(n423) );
  AOI21_X1 U397 ( .B1(n366), .B2(n423), .A(n365), .ZN(n346) );
  AOI22_X1 U398 ( .A1(n111), .A2(rs1_val_i[20]), .B1(n112), .B2(pc_i[20]), 
        .ZN(n345) );
  OAI21_X1 U399 ( .B1(n56), .B2(n346), .A(n345), .ZN(n599) );
  INV_X1 U400 ( .A(rs1_val_i[21]), .ZN(n425) );
  AOI21_X1 U401 ( .B1(n366), .B2(n425), .A(n365), .ZN(n348) );
  AOI22_X1 U402 ( .A1(n111), .A2(rs1_val_i[21]), .B1(n112), .B2(pc_i[21]), 
        .ZN(n347) );
  OAI21_X1 U403 ( .B1(n55), .B2(n348), .A(n347), .ZN(n598) );
  INV_X1 U404 ( .A(rs1_val_i[22]), .ZN(n427) );
  AOI21_X1 U405 ( .B1(n366), .B2(n427), .A(n365), .ZN(n350) );
  AOI22_X1 U406 ( .A1(n111), .A2(rs1_val_i[22]), .B1(n112), .B2(pc_i[22]), 
        .ZN(n349) );
  OAI21_X1 U407 ( .B1(n54), .B2(n350), .A(n349), .ZN(n597) );
  INV_X1 U408 ( .A(rs1_val_i[23]), .ZN(n429) );
  AOI21_X1 U409 ( .B1(n366), .B2(n429), .A(n365), .ZN(n352) );
  AOI22_X1 U410 ( .A1(n111), .A2(rs1_val_i[23]), .B1(n112), .B2(pc_i[23]), 
        .ZN(n351) );
  OAI21_X1 U411 ( .B1(n53), .B2(n352), .A(n351), .ZN(n596) );
  INV_X1 U412 ( .A(rs1_val_i[24]), .ZN(n431) );
  AOI21_X1 U413 ( .B1(n366), .B2(n431), .A(n365), .ZN(n354) );
  AOI22_X1 U414 ( .A1(n111), .A2(rs1_val_i[24]), .B1(n112), .B2(pc_i[24]), 
        .ZN(n353) );
  OAI21_X1 U415 ( .B1(n52), .B2(n354), .A(n353), .ZN(n595) );
  INV_X1 U416 ( .A(rs1_val_i[25]), .ZN(n433) );
  AOI21_X1 U417 ( .B1(n366), .B2(n433), .A(n365), .ZN(n356) );
  AOI22_X1 U418 ( .A1(n111), .A2(rs1_val_i[25]), .B1(n112), .B2(pc_i[25]), 
        .ZN(n355) );
  OAI21_X1 U419 ( .B1(n51), .B2(n356), .A(n355), .ZN(n594) );
  INV_X1 U420 ( .A(rs1_val_i[26]), .ZN(n435) );
  AOI21_X1 U421 ( .B1(n366), .B2(n435), .A(n365), .ZN(n358) );
  AOI22_X1 U422 ( .A1(n111), .A2(rs1_val_i[26]), .B1(n374), .B2(pc_i[26]), 
        .ZN(n357) );
  OAI21_X1 U423 ( .B1(n50), .B2(n358), .A(n357), .ZN(n593) );
  INV_X1 U424 ( .A(rs1_val_i[27]), .ZN(n437) );
  AOI21_X1 U425 ( .B1(n366), .B2(n437), .A(n365), .ZN(n360) );
  AOI22_X1 U426 ( .A1(n111), .A2(rs1_val_i[27]), .B1(n374), .B2(pc_i[27]), 
        .ZN(n359) );
  OAI21_X1 U427 ( .B1(n49), .B2(n360), .A(n359), .ZN(n592) );
  INV_X1 U428 ( .A(rs1_val_i[28]), .ZN(n439) );
  AOI21_X1 U429 ( .B1(n366), .B2(n439), .A(n110), .ZN(n362) );
  AOI22_X1 U430 ( .A1(n111), .A2(rs1_val_i[28]), .B1(n374), .B2(pc_i[28]), 
        .ZN(n361) );
  OAI21_X1 U431 ( .B1(n48), .B2(n362), .A(n361), .ZN(n591) );
  INV_X1 U432 ( .A(rs1_val_i[29]), .ZN(n441) );
  AOI21_X1 U433 ( .B1(n366), .B2(n441), .A(n365), .ZN(n364) );
  AOI22_X1 U434 ( .A1(n111), .A2(rs1_val_i[29]), .B1(n374), .B2(pc_i[29]), 
        .ZN(n363) );
  OAI21_X1 U435 ( .B1(n47), .B2(n364), .A(n363), .ZN(n590) );
  INV_X1 U436 ( .A(rs1_val_i[30]), .ZN(n444) );
  AOI21_X1 U437 ( .B1(n366), .B2(n444), .A(n110), .ZN(n369) );
  AOI22_X1 U438 ( .A1(n111), .A2(rs1_val_i[30]), .B1(n374), .B2(pc_i[30]), 
        .ZN(n368) );
  OAI21_X1 U439 ( .B1(n46), .B2(n369), .A(n368), .ZN(n589) );
  INV_X1 U440 ( .A(n449), .ZN(n372) );
  OAI21_X1 U441 ( .B1(n372), .B2(n371), .A(n370), .ZN(n373) );
  AOI22_X1 U442 ( .A1(n112), .A2(pc_i[31]), .B1(csr_mepc_o[31]), .B2(n373), 
        .ZN(n375) );
  OAI21_X1 U443 ( .B1(n376), .B2(n449), .A(n375), .ZN(n588) );
  OAI221_X1 U444 ( .B1(n447), .B2(n378), .C1(n447), .C2(n446), .A(csr_sr_q[4]), 
        .ZN(n377) );
  OAI21_X1 U445 ( .B1(n378), .B2(n450), .A(n377), .ZN(n587) );
  OAI221_X1 U446 ( .B1(n79), .B2(n446), .C1(n79), .C2(n382), .A(csr_sr_q[5]), 
        .ZN(n381) );
  OAI21_X1 U447 ( .B1(n445), .B2(n382), .A(n381), .ZN(n586) );
  OAI221_X1 U448 ( .B1(n79), .B2(n446), .C1(n79), .C2(n384), .A(csr_sr_q[6]), 
        .ZN(n383) );
  OAI21_X1 U449 ( .B1(n445), .B2(n384), .A(n383), .ZN(n585) );
  OAI21_X1 U450 ( .B1(n387), .B2(n386), .A(n385), .ZN(n404) );
  AOI21_X1 U451 ( .B1(n446), .B2(n393), .A(n404), .ZN(n392) );
  AOI21_X1 U452 ( .B1(csr_sr_q[3]), .B2(n389), .A(n388), .ZN(n390) );
  OAI222_X1 U453 ( .A1(n445), .A2(n393), .B1(n106), .B2(n392), .C1(n391), .C2(
        n390), .ZN(n584) );
  OAI221_X1 U454 ( .B1(n79), .B2(n446), .C1(n79), .C2(n395), .A(csr_sr_q[8]), 
        .ZN(n394) );
  OAI21_X1 U455 ( .B1(n445), .B2(n395), .A(n394), .ZN(n583) );
  OAI221_X1 U456 ( .B1(n79), .B2(n446), .C1(n79), .C2(n397), .A(csr_sr_q[9]), 
        .ZN(n396) );
  OAI21_X1 U457 ( .B1(n445), .B2(n397), .A(n396), .ZN(n582) );
  OAI221_X1 U458 ( .B1(n79), .B2(n446), .C1(n442), .C2(n399), .A(csr_sr_q[10]), 
        .ZN(n398) );
  OAI21_X1 U459 ( .B1(n445), .B2(n399), .A(n398), .ZN(n581) );
  NAND2_X1 U460 ( .A1(n401), .A2(n400), .ZN(n406) );
  OAI221_X1 U461 ( .B1(n404), .B2(n446), .C1(n404), .C2(n403), .A(csr_sr_q[11]), .ZN(n402) );
  OAI211_X1 U462 ( .C1(n445), .C2(n403), .A(n406), .B(n402), .ZN(n580) );
  OAI221_X1 U463 ( .B1(n404), .B2(n446), .C1(n404), .C2(n407), .A(csr_sr_q[12]), .ZN(n405) );
  OAI211_X1 U464 ( .C1(n445), .C2(n407), .A(n406), .B(n405), .ZN(n579) );
  OAI221_X1 U465 ( .B1(n79), .B2(n446), .C1(n442), .C2(n409), .A(csr_sr_q[13]), 
        .ZN(n408) );
  OAI21_X1 U466 ( .B1(n445), .B2(n409), .A(n408), .ZN(n578) );
  OAI221_X1 U467 ( .B1(n79), .B2(n446), .C1(n442), .C2(n411), .A(csr_sr_q[14]), 
        .ZN(n410) );
  OAI21_X1 U468 ( .B1(n445), .B2(n411), .A(n410), .ZN(n577) );
  OAI221_X1 U469 ( .B1(n79), .B2(n446), .C1(n79), .C2(n413), .A(csr_sr_q[15]), 
        .ZN(n412) );
  OAI21_X1 U470 ( .B1(n445), .B2(n413), .A(n412), .ZN(n576) );
  OAI221_X1 U471 ( .B1(n79), .B2(n446), .C1(n79), .C2(n415), .A(csr_sr_q[16]), 
        .ZN(n414) );
  OAI21_X1 U472 ( .B1(n445), .B2(n415), .A(n414), .ZN(n575) );
  OAI221_X1 U473 ( .B1(n79), .B2(n446), .C1(n79), .C2(n417), .A(csr_sr_q[17]), 
        .ZN(n416) );
  OAI21_X1 U474 ( .B1(n445), .B2(n417), .A(n416), .ZN(n574) );
  OAI221_X1 U475 ( .B1(n79), .B2(n446), .C1(n79), .C2(n419), .A(csr_sr_q[18]), 
        .ZN(n418) );
  OAI21_X1 U476 ( .B1(n445), .B2(n419), .A(n418), .ZN(n573) );
  OAI221_X1 U477 ( .B1(n79), .B2(n446), .C1(n79), .C2(n421), .A(csr_sr_q[19]), 
        .ZN(n420) );
  OAI21_X1 U478 ( .B1(n445), .B2(n421), .A(n420), .ZN(n572) );
  OAI221_X1 U479 ( .B1(n79), .B2(n446), .C1(n442), .C2(n423), .A(csr_sr_q[20]), 
        .ZN(n422) );
  OAI21_X1 U480 ( .B1(n445), .B2(n423), .A(n422), .ZN(n571) );
  OAI221_X1 U481 ( .B1(n79), .B2(n446), .C1(n79), .C2(n425), .A(csr_sr_q[21]), 
        .ZN(n424) );
  OAI21_X1 U482 ( .B1(n445), .B2(n425), .A(n424), .ZN(n570) );
  OAI221_X1 U483 ( .B1(n79), .B2(n446), .C1(n442), .C2(n427), .A(csr_sr_q[22]), 
        .ZN(n426) );
  OAI21_X1 U484 ( .B1(n445), .B2(n427), .A(n426), .ZN(n569) );
  OAI221_X1 U485 ( .B1(n79), .B2(n446), .C1(n79), .C2(n429), .A(csr_sr_q[23]), 
        .ZN(n428) );
  OAI21_X1 U486 ( .B1(n445), .B2(n429), .A(n428), .ZN(n568) );
  OAI221_X1 U487 ( .B1(n79), .B2(n446), .C1(n442), .C2(n431), .A(csr_sr_q[24]), 
        .ZN(n430) );
  OAI21_X1 U488 ( .B1(n445), .B2(n431), .A(n430), .ZN(n567) );
  OAI221_X1 U489 ( .B1(n79), .B2(n446), .C1(n442), .C2(n433), .A(csr_sr_q[25]), 
        .ZN(n432) );
  OAI21_X1 U490 ( .B1(n445), .B2(n433), .A(n432), .ZN(n566) );
  OAI221_X1 U491 ( .B1(n79), .B2(n446), .C1(n79), .C2(n435), .A(csr_sr_q[26]), 
        .ZN(n434) );
  OAI21_X1 U492 ( .B1(n445), .B2(n435), .A(n434), .ZN(n565) );
  OAI221_X1 U493 ( .B1(n79), .B2(n446), .C1(n442), .C2(n437), .A(csr_sr_q[27]), 
        .ZN(n436) );
  OAI21_X1 U494 ( .B1(n445), .B2(n437), .A(n436), .ZN(n564) );
  OAI221_X1 U495 ( .B1(n79), .B2(n446), .C1(n442), .C2(n439), .A(csr_sr_q[28]), 
        .ZN(n438) );
  OAI21_X1 U496 ( .B1(n445), .B2(n439), .A(n438), .ZN(n563) );
  OAI221_X1 U497 ( .B1(n79), .B2(n446), .C1(n442), .C2(n441), .A(csr_sr_q[29]), 
        .ZN(n440) );
  OAI21_X1 U498 ( .B1(n445), .B2(n441), .A(n440), .ZN(n562) );
  OAI221_X1 U499 ( .B1(n79), .B2(n446), .C1(n442), .C2(n444), .A(csr_sr_q[30]), 
        .ZN(n443) );
  OAI21_X1 U500 ( .B1(n445), .B2(n444), .A(n443), .ZN(n561) );
  OAI221_X1 U501 ( .B1(n447), .B2(n446), .C1(n447), .C2(n449), .A(csr_sr_q[31]), .ZN(n448) );
  OAI21_X1 U502 ( .B1(n450), .B2(n449), .A(n448), .ZN(n560) );
endmodule


module uriscv_muldiv ( clk_i, rst_i, valid_i, inst_mul_i, inst_mulh_i, 
        inst_mulhsu_i, inst_mulhu_i, inst_div_i, inst_divu_i, inst_rem_i, 
        inst_remu_i, operand_ra_i, operand_rb_i, stall_o, ready_o, result_o );
  input [31:0] operand_ra_i;
  input [31:0] operand_rb_i;
  output [31:0] result_o;
  input clk_i, rst_i, valid_i, inst_mul_i, inst_mulh_i, inst_mulhsu_i,
         inst_mulhu_i, inst_div_i, inst_divu_i, inst_rem_i, inst_remu_i;
  output stall_o, ready_o;
  wire   mulhi_sel_q, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66,
         N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80,
         N81, N82, N83, N84, N85, N86, N88, N89, mul_busy_q, div_busy_q,
         div_inst_q, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200,
         N575, C22_DATA3_1, C22_DATA3_2, C22_DATA3_3, C22_DATA3_4, C22_DATA3_5,
         C22_DATA3_6, C22_DATA3_7, C22_DATA3_8, C22_DATA3_9, C22_DATA3_10,
         C22_DATA3_11, C22_DATA3_12, C22_DATA3_13, C22_DATA3_14, C22_DATA3_15,
         C22_DATA3_16, C22_DATA3_17, C22_DATA3_18, C22_DATA3_19, C22_DATA3_20,
         C22_DATA3_21, C22_DATA3_22, C22_DATA3_23, C22_DATA3_24, C22_DATA3_25,
         C22_DATA3_26, C22_DATA3_27, C22_DATA3_28, C22_DATA3_29, C22_DATA3_30,
         C21_DATA3_0, C21_DATA3_1, C21_DATA3_2, C21_DATA3_3, C21_DATA3_4,
         C21_DATA3_5, C21_DATA3_6, C21_DATA3_7, C21_DATA3_8, C21_DATA3_9,
         C21_DATA3_10, C21_DATA3_11, C21_DATA3_12, C21_DATA3_13, C21_DATA3_14,
         C21_DATA3_15, C21_DATA3_16, C21_DATA3_17, C21_DATA3_18, C21_DATA3_19,
         C21_DATA3_20, C21_DATA3_21, C21_DATA3_22, C21_DATA3_23, C21_DATA3_24,
         C21_DATA3_25, C21_DATA3_26, C21_DATA3_27, C21_DATA3_28, C21_DATA3_29,
         C21_DATA3_30, n6400, n7100, n7200, n7300, n7400, n7500, n7600, n7700,
         n7800, n7900, n8000, n8100, n8200, n8300, n8400, n8500, n8600, n87,
         n8800, n8900, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n290, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n386, n402, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n5750, n576, n577,
         n578, C1_Z_31, C1_Z_30, C1_Z_29, C1_Z_28, C1_Z_27, C1_Z_26, C1_Z_25,
         C1_Z_24, C1_Z_23, C1_Z_22, C1_Z_21, C1_Z_20, C1_Z_19, C1_Z_18,
         C1_Z_17, C1_Z_16, C1_Z_15, C1_Z_14, C1_Z_13, C1_Z_12, C1_Z_11,
         C1_Z_10, C1_Z_9, C1_Z_8, C1_Z_7, C1_Z_6, C1_Z_5, C1_Z_4, C1_Z_3,
         C1_Z_2, C1_Z_1, C1_Z_0, sub_x_9_n30, sub_x_9_n29, sub_x_9_n28,
         sub_x_9_n27, sub_x_9_n26, sub_x_9_n25, sub_x_9_n24, sub_x_9_n23,
         sub_x_9_n22, sub_x_9_n21, sub_x_9_n20, sub_x_9_n19, sub_x_9_n18,
         sub_x_9_n17, sub_x_9_n16, sub_x_9_n15, sub_x_9_n14, sub_x_9_n13,
         sub_x_9_n12, sub_x_9_n11, sub_x_9_n10, sub_x_9_n9, sub_x_9_n8,
         sub_x_9_n7, sub_x_9_n6, sub_x_9_n5, sub_x_9_n4, sub_x_9_n3,
         sub_x_9_n2, sub_x_9_n1, DP_OP_63J3_127_9516_n30,
         DP_OP_63J3_127_9516_n29, DP_OP_63J3_127_9516_n28,
         DP_OP_63J3_127_9516_n27, DP_OP_63J3_127_9516_n26,
         DP_OP_63J3_127_9516_n25, DP_OP_63J3_127_9516_n24,
         DP_OP_63J3_127_9516_n23, DP_OP_63J3_127_9516_n22,
         DP_OP_63J3_127_9516_n21, DP_OP_63J3_127_9516_n20,
         DP_OP_63J3_127_9516_n19, DP_OP_63J3_127_9516_n18,
         DP_OP_63J3_127_9516_n17, DP_OP_63J3_127_9516_n16,
         DP_OP_63J3_127_9516_n15, DP_OP_63J3_127_9516_n14,
         DP_OP_63J3_127_9516_n13, DP_OP_63J3_127_9516_n12,
         DP_OP_63J3_127_9516_n11, DP_OP_63J3_127_9516_n10,
         DP_OP_63J3_127_9516_n9, DP_OP_63J3_127_9516_n8,
         DP_OP_63J3_127_9516_n7, DP_OP_63J3_127_9516_n6,
         DP_OP_63J3_127_9516_n5, DP_OP_63J3_127_9516_n4,
         DP_OP_63J3_127_9516_n3, DP_OP_63J3_127_9516_n2,
         DP_OP_63J3_127_9516_n1, mult_x_6_n1483, mult_x_6_n1482,
         mult_x_6_n1481, mult_x_6_n1480, mult_x_6_n1479, mult_x_6_n1478,
         mult_x_6_n1477, mult_x_6_n1476, mult_x_6_n1475, mult_x_6_n1474,
         mult_x_6_n1473, mult_x_6_n1472, mult_x_6_n1471, mult_x_6_n1470,
         mult_x_6_n1469, mult_x_6_n1468, mult_x_6_n1467, mult_x_6_n1466,
         mult_x_6_n1465, mult_x_6_n1464, mult_x_6_n1463, mult_x_6_n1462,
         mult_x_6_n1461, mult_x_6_n1460, mult_x_6_n1459, mult_x_6_n1458,
         mult_x_6_n1457, mult_x_6_n1456, mult_x_6_n1455, mult_x_6_n1454,
         mult_x_6_n1453, mult_x_6_n1452, mult_x_6_n1451, mult_x_6_n1450,
         mult_x_6_n1447, mult_x_6_n1445, mult_x_6_n1444, mult_x_6_n1443,
         mult_x_6_n1442, mult_x_6_n1441, mult_x_6_n1440, mult_x_6_n1439,
         mult_x_6_n1437, mult_x_6_n1436, mult_x_6_n1435, mult_x_6_n1434,
         mult_x_6_n1433, mult_x_6_n1432, mult_x_6_n1431, mult_x_6_n1430,
         mult_x_6_n1429, mult_x_6_n1428, mult_x_6_n1427, mult_x_6_n1426,
         mult_x_6_n1425, mult_x_6_n1424, mult_x_6_n1423, mult_x_6_n1422,
         mult_x_6_n1421, mult_x_6_n1420, mult_x_6_n1419, mult_x_6_n1418,
         mult_x_6_n1417, mult_x_6_n1416, mult_x_6_n1415, mult_x_6_n1414,
         mult_x_6_n1413, mult_x_6_n1411, mult_x_6_n1410, mult_x_6_n1409,
         mult_x_6_n1408, mult_x_6_n1407, mult_x_6_n1406, mult_x_6_n1405,
         mult_x_6_n1404, mult_x_6_n1403, mult_x_6_n1402, mult_x_6_n1401,
         mult_x_6_n1400, mult_x_6_n1399, mult_x_6_n1398, mult_x_6_n1397,
         mult_x_6_n1396, mult_x_6_n1395, mult_x_6_n1394, mult_x_6_n1393,
         mult_x_6_n1392, mult_x_6_n1391, mult_x_6_n1390, mult_x_6_n1389,
         mult_x_6_n1388, mult_x_6_n1387, mult_x_6_n1386, mult_x_6_n1385,
         mult_x_6_n1384, mult_x_6_n1383, mult_x_6_n1382, mult_x_6_n1381,
         mult_x_6_n1380, mult_x_6_n1379, mult_x_6_n1376, mult_x_6_n1375,
         mult_x_6_n1374, mult_x_6_n1373, mult_x_6_n1372, mult_x_6_n1371,
         mult_x_6_n1370, mult_x_6_n1369, mult_x_6_n1368, mult_x_6_n1367,
         mult_x_6_n1366, mult_x_6_n1365, mult_x_6_n1364, mult_x_6_n1363,
         mult_x_6_n1362, mult_x_6_n1361, mult_x_6_n1360, mult_x_6_n1359,
         mult_x_6_n1358, mult_x_6_n1357, mult_x_6_n1356, mult_x_6_n1355,
         mult_x_6_n1354, mult_x_6_n1353, mult_x_6_n1352, mult_x_6_n1351,
         mult_x_6_n1350, mult_x_6_n1349, mult_x_6_n1348, mult_x_6_n1347,
         mult_x_6_n1346, mult_x_6_n1345, mult_x_6_n1344, mult_x_6_n1341,
         mult_x_6_n1340, mult_x_6_n1339, mult_x_6_n1338, mult_x_6_n1337,
         mult_x_6_n1336, mult_x_6_n1335, mult_x_6_n1334, mult_x_6_n1333,
         mult_x_6_n1332, mult_x_6_n1331, mult_x_6_n1330, mult_x_6_n1329,
         mult_x_6_n1328, mult_x_6_n1327, mult_x_6_n1326, mult_x_6_n1325,
         mult_x_6_n1324, mult_x_6_n1323, mult_x_6_n1322, mult_x_6_n1321,
         mult_x_6_n1320, mult_x_6_n1319, mult_x_6_n1318, mult_x_6_n1317,
         mult_x_6_n1316, mult_x_6_n1315, mult_x_6_n1314, mult_x_6_n1313,
         mult_x_6_n1312, mult_x_6_n1311, mult_x_6_n1310, mult_x_6_n1309,
         mult_x_6_n1306, mult_x_6_n1305, mult_x_6_n1304, mult_x_6_n1303,
         mult_x_6_n1302, mult_x_6_n1301, mult_x_6_n1300, mult_x_6_n1299,
         mult_x_6_n1298, mult_x_6_n1297, mult_x_6_n1296, mult_x_6_n1295,
         mult_x_6_n1294, mult_x_6_n1293, mult_x_6_n1292, mult_x_6_n1291,
         mult_x_6_n1290, mult_x_6_n1289, mult_x_6_n1288, mult_x_6_n1287,
         mult_x_6_n1286, mult_x_6_n1285, mult_x_6_n1284, mult_x_6_n1283,
         mult_x_6_n1282, mult_x_6_n1281, mult_x_6_n1280, mult_x_6_n1279,
         mult_x_6_n1278, mult_x_6_n1277, mult_x_6_n1276, mult_x_6_n1275,
         mult_x_6_n1274, mult_x_6_n1273, mult_x_6_n1272, mult_x_6_n1271,
         mult_x_6_n1270, mult_x_6_n1269, mult_x_6_n1268, mult_x_6_n1267,
         mult_x_6_n1266, mult_x_6_n1265, mult_x_6_n1264, mult_x_6_n1263,
         mult_x_6_n1262, mult_x_6_n1261, mult_x_6_n1260, mult_x_6_n1259,
         mult_x_6_n1258, mult_x_6_n1257, mult_x_6_n1256, mult_x_6_n1255,
         mult_x_6_n1254, mult_x_6_n1253, mult_x_6_n1252, mult_x_6_n1251,
         mult_x_6_n1250, mult_x_6_n1249, mult_x_6_n1248, mult_x_6_n1247,
         mult_x_6_n1246, mult_x_6_n1245, mult_x_6_n1244, mult_x_6_n1243,
         mult_x_6_n1242, mult_x_6_n1241, mult_x_6_n1240, mult_x_6_n1239,
         mult_x_6_n1238, mult_x_6_n1237, mult_x_6_n1236, mult_x_6_n1235,
         mult_x_6_n1234, mult_x_6_n1233, mult_x_6_n1232, mult_x_6_n1231,
         mult_x_6_n1230, mult_x_6_n1229, mult_x_6_n1228, mult_x_6_n1227,
         mult_x_6_n1226, mult_x_6_n1225, mult_x_6_n1224, mult_x_6_n1223,
         mult_x_6_n1222, mult_x_6_n1221, mult_x_6_n1220, mult_x_6_n1219,
         mult_x_6_n1218, mult_x_6_n1217, mult_x_6_n1216, mult_x_6_n1215,
         mult_x_6_n1214, mult_x_6_n1213, mult_x_6_n1212, mult_x_6_n1211,
         mult_x_6_n1210, mult_x_6_n1209, mult_x_6_n1208, mult_x_6_n1207,
         mult_x_6_n1206, mult_x_6_n1205, mult_x_6_n1204, mult_x_6_n1203,
         mult_x_6_n1202, mult_x_6_n1201, mult_x_6_n1200, mult_x_6_n1199,
         mult_x_6_n1198, mult_x_6_n1197, mult_x_6_n1196, mult_x_6_n1195,
         mult_x_6_n1194, mult_x_6_n1193, mult_x_6_n1192, mult_x_6_n1191,
         mult_x_6_n1190, mult_x_6_n1189, mult_x_6_n1188, mult_x_6_n1187,
         mult_x_6_n1186, mult_x_6_n1185, mult_x_6_n1184, mult_x_6_n1183,
         mult_x_6_n1182, mult_x_6_n1181, mult_x_6_n1180, mult_x_6_n1179,
         mult_x_6_n1178, mult_x_6_n1177, mult_x_6_n1176, mult_x_6_n1175,
         mult_x_6_n1174, mult_x_6_n1173, mult_x_6_n1172, mult_x_6_n1171,
         mult_x_6_n1170, mult_x_6_n1169, mult_x_6_n1168, mult_x_6_n1167,
         mult_x_6_n1166, mult_x_6_n1165, mult_x_6_n1164, mult_x_6_n1163,
         mult_x_6_n1162, mult_x_6_n1161, mult_x_6_n1160, mult_x_6_n1159,
         mult_x_6_n1158, mult_x_6_n1157, mult_x_6_n1156, mult_x_6_n1155,
         mult_x_6_n1154, mult_x_6_n1153, mult_x_6_n1152, mult_x_6_n1151,
         mult_x_6_n1150, mult_x_6_n1149, mult_x_6_n1148, mult_x_6_n1147,
         mult_x_6_n1146, mult_x_6_n1145, mult_x_6_n1144, mult_x_6_n1143,
         mult_x_6_n1142, mult_x_6_n1141, mult_x_6_n1140, mult_x_6_n1139,
         mult_x_6_n1138, mult_x_6_n1137, mult_x_6_n1136, mult_x_6_n1135,
         mult_x_6_n1134, mult_x_6_n1133, mult_x_6_n1132, mult_x_6_n1131,
         mult_x_6_n1130, mult_x_6_n1129, mult_x_6_n1128, mult_x_6_n1127,
         mult_x_6_n1126, mult_x_6_n1125, mult_x_6_n1124, mult_x_6_n1123,
         mult_x_6_n1122, mult_x_6_n1121, mult_x_6_n1120, mult_x_6_n1119,
         mult_x_6_n1118, mult_x_6_n1117, mult_x_6_n1116, mult_x_6_n1115,
         mult_x_6_n1114, mult_x_6_n1113, mult_x_6_n1112, mult_x_6_n1111,
         mult_x_6_n1110, mult_x_6_n1109, mult_x_6_n1108, mult_x_6_n1107,
         mult_x_6_n1106, mult_x_6_n1103, mult_x_6_n1102, mult_x_6_n1101,
         mult_x_6_n1100, mult_x_6_n1098, mult_x_6_n1097, mult_x_6_n1096,
         mult_x_6_n1095, mult_x_6_n1094, mult_x_6_n1093, mult_x_6_n1092,
         mult_x_6_n1091, mult_x_6_n1090, mult_x_6_n1089, mult_x_6_n1088,
         mult_x_6_n1087, mult_x_6_n1086, mult_x_6_n1085, mult_x_6_n1084,
         mult_x_6_n1083, mult_x_6_n1082, mult_x_6_n1081, mult_x_6_n1080,
         mult_x_6_n1079, mult_x_6_n1078, mult_x_6_n1077, mult_x_6_n1076,
         mult_x_6_n1075, mult_x_6_n1074, mult_x_6_n1073, mult_x_6_n1072,
         mult_x_6_n1071, mult_x_6_n1070, mult_x_6_n1069, mult_x_6_n1067,
         mult_x_6_n1064, mult_x_6_n1063, mult_x_6_n1059, mult_x_6_n1058,
         mult_x_6_n1057, mult_x_6_n1056, mult_x_6_n1055, mult_x_6_n1054,
         mult_x_6_n1053, mult_x_6_n1051, mult_x_6_n1050, mult_x_6_n1049,
         mult_x_6_n1047, mult_x_6_n1046, mult_x_6_n1044, mult_x_6_n1042,
         mult_x_6_n1041, mult_x_6_n1040, mult_x_6_n995, mult_x_6_n994,
         mult_x_6_n993, mult_x_6_n991, mult_x_6_n989, mult_x_6_n988,
         mult_x_6_n987, mult_x_6_n986, mult_x_6_n985, mult_x_6_n984,
         mult_x_6_n983, mult_x_6_n982, mult_x_6_n981, mult_x_6_n980,
         mult_x_6_n979, mult_x_6_n978, mult_x_6_n977, mult_x_6_n976,
         mult_x_6_n975, mult_x_6_n974, mult_x_6_n973, mult_x_6_n972,
         mult_x_6_n971, mult_x_6_n970, mult_x_6_n969, mult_x_6_n967,
         mult_x_6_n966, mult_x_6_n965, mult_x_6_n964, mult_x_6_n963,
         mult_x_6_n962, mult_x_6_n961, mult_x_6_n960, mult_x_6_n959,
         mult_x_6_n958, mult_x_6_n957, mult_x_6_n956, mult_x_6_n955,
         mult_x_6_n954, mult_x_6_n953, mult_x_6_n951, mult_x_6_n950,
         mult_x_6_n949, mult_x_6_n948, mult_x_6_n947, mult_x_6_n946,
         mult_x_6_n945, mult_x_6_n943, mult_x_6_n942, mult_x_6_n941,
         mult_x_6_n940, mult_x_6_n939, mult_x_6_n938, mult_x_6_n937,
         mult_x_6_n936, mult_x_6_n935, mult_x_6_n934, mult_x_6_n933,
         mult_x_6_n932, mult_x_6_n931, mult_x_6_n930, mult_x_6_n929,
         mult_x_6_n928, mult_x_6_n927, mult_x_6_n926, mult_x_6_n925,
         mult_x_6_n924, mult_x_6_n923, mult_x_6_n922, mult_x_6_n921,
         mult_x_6_n920, mult_x_6_n919, mult_x_6_n918, mult_x_6_n917,
         mult_x_6_n916, mult_x_6_n915, mult_x_6_n914, mult_x_6_n913,
         mult_x_6_n912, mult_x_6_n911, mult_x_6_n910, mult_x_6_n909,
         mult_x_6_n908, mult_x_6_n907, mult_x_6_n906, mult_x_6_n905,
         mult_x_6_n904, mult_x_6_n903, mult_x_6_n902, mult_x_6_n901,
         mult_x_6_n900, mult_x_6_n899, mult_x_6_n897, mult_x_6_n896,
         mult_x_6_n895, mult_x_6_n894, mult_x_6_n893, mult_x_6_n892,
         mult_x_6_n891, mult_x_6_n890, mult_x_6_n889, mult_x_6_n888,
         mult_x_6_n887, mult_x_6_n886, mult_x_6_n885, mult_x_6_n884,
         mult_x_6_n883, mult_x_6_n882, mult_x_6_n881, mult_x_6_n880,
         mult_x_6_n879, mult_x_6_n878, mult_x_6_n877, mult_x_6_n876,
         mult_x_6_n875, mult_x_6_n874, mult_x_6_n873, mult_x_6_n872,
         mult_x_6_n871, mult_x_6_n870, mult_x_6_n869, mult_x_6_n868,
         mult_x_6_n867, mult_x_6_n866, mult_x_6_n865, mult_x_6_n864,
         mult_x_6_n863, mult_x_6_n862, mult_x_6_n861, mult_x_6_n860,
         mult_x_6_n859, mult_x_6_n858, mult_x_6_n857, mult_x_6_n856,
         mult_x_6_n855, mult_x_6_n854, mult_x_6_n853, mult_x_6_n852,
         mult_x_6_n851, mult_x_6_n850, mult_x_6_n849, mult_x_6_n848,
         mult_x_6_n847, mult_x_6_n846, mult_x_6_n845, mult_x_6_n844,
         mult_x_6_n843, mult_x_6_n842, mult_x_6_n841, mult_x_6_n840,
         mult_x_6_n839, mult_x_6_n838, mult_x_6_n837, mult_x_6_n836,
         mult_x_6_n835, mult_x_6_n833, mult_x_6_n832, mult_x_6_n831,
         mult_x_6_n830, mult_x_6_n829, mult_x_6_n828, mult_x_6_n827,
         mult_x_6_n826, mult_x_6_n825, mult_x_6_n824, mult_x_6_n823,
         mult_x_6_n822, mult_x_6_n821, mult_x_6_n820, mult_x_6_n819,
         mult_x_6_n817, mult_x_6_n816, mult_x_6_n815, mult_x_6_n813,
         mult_x_6_n812, mult_x_6_n811, mult_x_6_n810, mult_x_6_n809,
         mult_x_6_n808, mult_x_6_n807, mult_x_6_n806, mult_x_6_n805,
         mult_x_6_n804, mult_x_6_n803, mult_x_6_n802, mult_x_6_n801,
         mult_x_6_n799, mult_x_6_n797, mult_x_6_n795, mult_x_6_n794,
         mult_x_6_n793, mult_x_6_n792, mult_x_6_n791, mult_x_6_n790,
         mult_x_6_n789, mult_x_6_n788, mult_x_6_n787, mult_x_6_n785,
         mult_x_6_n784, mult_x_6_n783, mult_x_6_n782, mult_x_6_n781,
         mult_x_6_n779, mult_x_6_n778, mult_x_6_n777, mult_x_6_n776,
         mult_x_6_n775, mult_x_6_n774, mult_x_6_n773, mult_x_6_n772,
         mult_x_6_n771, mult_x_6_n770, mult_x_6_n769, mult_x_6_n768,
         mult_x_6_n767, mult_x_6_n766, mult_x_6_n765, mult_x_6_n764,
         mult_x_6_n763, mult_x_6_n762, mult_x_6_n761, mult_x_6_n760,
         mult_x_6_n759, mult_x_6_n758, mult_x_6_n757, mult_x_6_n756,
         mult_x_6_n755, mult_x_6_n754, mult_x_6_n753, mult_x_6_n752,
         mult_x_6_n751, mult_x_6_n750, mult_x_6_n749, mult_x_6_n747,
         mult_x_6_n746, mult_x_6_n745, mult_x_6_n744, mult_x_6_n743,
         mult_x_6_n742, mult_x_6_n741, mult_x_6_n740, mult_x_6_n739,
         mult_x_6_n738, mult_x_6_n737, mult_x_6_n736, mult_x_6_n735,
         mult_x_6_n734, mult_x_6_n733, mult_x_6_n732, mult_x_6_n731,
         mult_x_6_n730, mult_x_6_n729, mult_x_6_n728, mult_x_6_n727,
         mult_x_6_n726, mult_x_6_n725, mult_x_6_n724, mult_x_6_n723,
         mult_x_6_n722, mult_x_6_n721, mult_x_6_n720, mult_x_6_n719,
         mult_x_6_n718, mult_x_6_n717, mult_x_6_n716, mult_x_6_n715,
         mult_x_6_n714, mult_x_6_n713, mult_x_6_n712, mult_x_6_n711,
         mult_x_6_n710, mult_x_6_n709, mult_x_6_n708, mult_x_6_n707,
         mult_x_6_n706, mult_x_6_n705, mult_x_6_n704, mult_x_6_n703,
         mult_x_6_n702, mult_x_6_n701, mult_x_6_n700, mult_x_6_n699,
         mult_x_6_n698, mult_x_6_n697, mult_x_6_n696, mult_x_6_n695,
         mult_x_6_n694, mult_x_6_n693, mult_x_6_n692, mult_x_6_n691,
         mult_x_6_n689, mult_x_6_n688, mult_x_6_n687, mult_x_6_n686,
         mult_x_6_n685, mult_x_6_n684, mult_x_6_n683, mult_x_6_n682,
         mult_x_6_n681, mult_x_6_n680, mult_x_6_n679, mult_x_6_n678,
         mult_x_6_n677, mult_x_6_n676, mult_x_6_n675, mult_x_6_n674,
         mult_x_6_n673, mult_x_6_n672, mult_x_6_n671, mult_x_6_n670,
         mult_x_6_n669, mult_x_6_n667, mult_x_6_n666, mult_x_6_n665,
         mult_x_6_n664, mult_x_6_n663, mult_x_6_n662, mult_x_6_n661,
         mult_x_6_n660, mult_x_6_n659, mult_x_6_n658, mult_x_6_n657,
         mult_x_6_n656, mult_x_6_n655, mult_x_6_n654, mult_x_6_n653,
         mult_x_6_n652, mult_x_6_n651, mult_x_6_n650, mult_x_6_n649,
         mult_x_6_n648, mult_x_6_n647, mult_x_6_n646, mult_x_6_n645,
         mult_x_6_n644, mult_x_6_n643, mult_x_6_n642, mult_x_6_n641,
         mult_x_6_n640, mult_x_6_n639, mult_x_6_n638, mult_x_6_n637,
         mult_x_6_n636, mult_x_6_n635, mult_x_6_n634, mult_x_6_n633,
         mult_x_6_n632, mult_x_6_n631, mult_x_6_n630, mult_x_6_n629,
         mult_x_6_n628, mult_x_6_n627, mult_x_6_n625, mult_x_6_n624,
         mult_x_6_n623, mult_x_6_n622, mult_x_6_n621, mult_x_6_n620,
         mult_x_6_n619, mult_x_6_n618, mult_x_6_n617, mult_x_6_n616,
         mult_x_6_n615, mult_x_6_n614, mult_x_6_n613, mult_x_6_n612,
         mult_x_6_n611, mult_x_6_n610, mult_x_6_n609, mult_x_6_n608,
         mult_x_6_n606, mult_x_6_n605, mult_x_6_n604, mult_x_6_n603,
         mult_x_6_n602, mult_x_6_n601, mult_x_6_n600, mult_x_6_n599,
         mult_x_6_n598, mult_x_6_n597, mult_x_6_n596, mult_x_6_n595,
         mult_x_6_n594, mult_x_6_n593, mult_x_6_n592, mult_x_6_n591,
         mult_x_6_n590, mult_x_6_n589, mult_x_6_n588, mult_x_6_n587,
         mult_x_6_n586, mult_x_6_n585, mult_x_6_n584, mult_x_6_n583,
         mult_x_6_n582, mult_x_6_n581, mult_x_6_n580, mult_x_6_n579,
         mult_x_6_n578, mult_x_6_n577, mult_x_6_n576, mult_x_6_n575,
         mult_x_6_n574, mult_x_6_n573, mult_x_6_n572, mult_x_6_n571,
         mult_x_6_n570, mult_x_6_n568, mult_x_6_n567, mult_x_6_n566,
         mult_x_6_n565, mult_x_6_n564, mult_x_6_n563, mult_x_6_n562,
         mult_x_6_n561, mult_x_6_n560, mult_x_6_n559, mult_x_6_n558,
         mult_x_6_n557, mult_x_6_n556, mult_x_6_n555, mult_x_6_n554,
         mult_x_6_n553, mult_x_6_n551, mult_x_6_n550, mult_x_6_n549,
         mult_x_6_n548, mult_x_6_n547, mult_x_6_n546, mult_x_6_n545,
         mult_x_6_n544, mult_x_6_n543, mult_x_6_n542, mult_x_6_n541,
         mult_x_6_n540, mult_x_6_n539, mult_x_6_n538, mult_x_6_n537,
         mult_x_6_n536, mult_x_6_n535, mult_x_6_n534, mult_x_6_n533,
         mult_x_6_n532, mult_x_6_n531, mult_x_6_n530, mult_x_6_n529,
         mult_x_6_n528, mult_x_6_n527, mult_x_6_n526, mult_x_6_n525,
         mult_x_6_n524, mult_x_6_n523, mult_x_6_n522, mult_x_6_n521,
         mult_x_6_n520, mult_x_6_n518, mult_x_6_n517, mult_x_6_n516,
         mult_x_6_n515, mult_x_6_n514, mult_x_6_n513, mult_x_6_n512,
         mult_x_6_n511, mult_x_6_n510, mult_x_6_n509, mult_x_6_n508,
         mult_x_6_n507, mult_x_6_n506, mult_x_6_n505, mult_x_6_n503,
         mult_x_6_n502, mult_x_6_n501, mult_x_6_n500, mult_x_6_n499,
         mult_x_6_n498, mult_x_6_n497, mult_x_6_n496, mult_x_6_n495,
         mult_x_6_n494, mult_x_6_n493, mult_x_6_n492, mult_x_6_n491,
         mult_x_6_n490, mult_x_6_n489, mult_x_6_n488, mult_x_6_n487,
         mult_x_6_n486, mult_x_6_n485, mult_x_6_n484, mult_x_6_n483,
         mult_x_6_n482, mult_x_6_n481, mult_x_6_n480, mult_x_6_n479,
         mult_x_6_n478, mult_x_6_n477, mult_x_6_n476, mult_x_6_n475,
         mult_x_6_n473, mult_x_6_n472, mult_x_6_n471, mult_x_6_n470,
         mult_x_6_n469, mult_x_6_n468, mult_x_6_n467, mult_x_6_n466,
         mult_x_6_n465, mult_x_6_n464, mult_x_6_n463, mult_x_6_n462,
         mult_x_6_n460, mult_x_6_n459, mult_x_6_n458, mult_x_6_n457,
         mult_x_6_n456, mult_x_6_n455, mult_x_6_n454, mult_x_6_n453,
         mult_x_6_n452, mult_x_6_n451, mult_x_6_n450, mult_x_6_n449,
         mult_x_6_n448, mult_x_6_n447, mult_x_6_n446, mult_x_6_n445,
         mult_x_6_n444, mult_x_6_n443, mult_x_6_n442, mult_x_6_n441,
         mult_x_6_n440, mult_x_6_n439, mult_x_6_n438, mult_x_6_n437,
         mult_x_6_n435, mult_x_6_n434, mult_x_6_n433, mult_x_6_n432,
         mult_x_6_n431, mult_x_6_n430, mult_x_6_n429, mult_x_6_n428,
         mult_x_6_n427, mult_x_6_n426, mult_x_6_n424, mult_x_6_n423,
         mult_x_6_n422, mult_x_6_n421, mult_x_6_n420, mult_x_6_n419,
         mult_x_6_n418, mult_x_6_n417, mult_x_6_n416, mult_x_6_n415,
         mult_x_6_n414, mult_x_6_n413, mult_x_6_n412, mult_x_6_n411,
         mult_x_6_n410, mult_x_6_n409, mult_x_6_n408, mult_x_6_n407,
         mult_x_6_n406, mult_x_6_n405, mult_x_6_n404, mult_x_6_n402,
         mult_x_6_n401, mult_x_6_n400, mult_x_6_n399, mult_x_6_n398,
         mult_x_6_n397, mult_x_6_n396, mult_x_6_n395, mult_x_6_n393,
         mult_x_6_n392, mult_x_6_n391, mult_x_6_n390, mult_x_6_n389,
         mult_x_6_n388, mult_x_6_n387, mult_x_6_n386, mult_x_6_n385,
         mult_x_6_n384, mult_x_6_n383, mult_x_6_n382, mult_x_6_n381,
         mult_x_6_n380, mult_x_6_n379, mult_x_6_n378, mult_x_6_n376,
         mult_x_6_n375, mult_x_6_n374, mult_x_6_n373, mult_x_6_n372,
         mult_x_6_n371, mult_x_6_n369, mult_x_6_n368, mult_x_6_n367,
         mult_x_6_n366, mult_x_6_n365, mult_x_6_n364, mult_x_6_n363,
         mult_x_6_n362, mult_x_6_n361, mult_x_6_n360, mult_x_6_n359,
         mult_x_6_n358, mult_x_6_n357, mult_x_6_n355, mult_x_6_n354,
         mult_x_6_n353, mult_x_6_n352, mult_x_6_n350, mult_x_6_n349,
         mult_x_6_n348, mult_x_6_n347, mult_x_6_n346, mult_x_6_n345,
         mult_x_6_n344, mult_x_6_n343, mult_x_6_n341, mult_x_6_n340,
         mult_x_6_n338, mult_x_6_n337, mult_x_6_n336, mult_x_6_n335,
         mult_x_6_n334, mult_x_6_n333, mult_x_6_n330, mult_x_6_n329,
         mult_x_6_n328, mult_x_6_n327, mult_x_6_n326, mult_x_6_n325,
         mult_x_6_n324, mult_x_6_n323, mult_x_6_n321, mult_x_6_n318,
         mult_x_6_n316, mult_x_6_n314, mult_x_6_n313, mult_x_6_n312,
         mult_x_6_n309, mult_x_6_n308, mult_x_6_n307, mult_x_6_n306,
         mult_x_6_n304, mult_x_6_n301, mult_x_6_n300, mult_x_6_n299,
         mult_x_6_n297, mult_x_6_n295, mult_x_6_n294, mult_x_6_n292,
         mult_x_6_n286, mult_x_6_n285, mult_x_6_n283, mult_x_6_n282,
         mult_x_6_n281, mult_x_6_n280, mult_x_6_n278, mult_x_6_n277,
         mult_x_6_n276, mult_x_6_n275, mult_x_6_n273, mult_x_6_n270,
         DP_OP_56J3_124_887_n132, DP_OP_56J3_124_887_n131,
         DP_OP_56J3_124_887_n130, DP_OP_56J3_124_887_n129,
         DP_OP_56J3_124_887_n128, DP_OP_56J3_124_887_n127,
         DP_OP_56J3_124_887_n126, DP_OP_56J3_124_887_n125,
         DP_OP_56J3_124_887_n124, DP_OP_56J3_124_887_n123,
         DP_OP_56J3_124_887_n122, DP_OP_56J3_124_887_n121,
         DP_OP_56J3_124_887_n120, DP_OP_56J3_124_887_n119,
         DP_OP_56J3_124_887_n118, DP_OP_56J3_124_887_n117,
         DP_OP_56J3_124_887_n116, DP_OP_56J3_124_887_n115,
         DP_OP_56J3_124_887_n114, DP_OP_56J3_124_887_n113,
         DP_OP_56J3_124_887_n112, DP_OP_56J3_124_887_n111,
         DP_OP_56J3_124_887_n110, DP_OP_56J3_124_887_n109,
         DP_OP_56J3_124_887_n108, DP_OP_56J3_124_887_n107,
         DP_OP_56J3_124_887_n106, DP_OP_56J3_124_887_n105,
         DP_OP_56J3_124_887_n104, DP_OP_56J3_124_887_n103,
         DP_OP_56J3_124_887_n102, DP_OP_56J3_124_887_n32,
         DP_OP_56J3_124_887_n31, DP_OP_56J3_124_887_n30,
         DP_OP_56J3_124_887_n29, DP_OP_56J3_124_887_n28,
         DP_OP_56J3_124_887_n27, DP_OP_56J3_124_887_n26,
         DP_OP_56J3_124_887_n25, DP_OP_56J3_124_887_n24,
         DP_OP_56J3_124_887_n23, DP_OP_56J3_124_887_n22,
         DP_OP_56J3_124_887_n21, DP_OP_56J3_124_887_n20,
         DP_OP_56J3_124_887_n19, DP_OP_56J3_124_887_n18,
         DP_OP_56J3_124_887_n17, DP_OP_56J3_124_887_n16,
         DP_OP_56J3_124_887_n15, DP_OP_56J3_124_887_n14,
         DP_OP_56J3_124_887_n13, DP_OP_56J3_124_887_n12,
         DP_OP_56J3_124_887_n11, DP_OP_56J3_124_887_n10, DP_OP_56J3_124_887_n9,
         DP_OP_56J3_124_887_n8, DP_OP_56J3_124_887_n7, DP_OP_56J3_124_887_n6,
         DP_OP_56J3_124_887_n5, DP_OP_56J3_124_887_n4, DP_OP_56J3_124_887_n3,
         DP_OP_56J3_124_887_n2, DP_OP_56J3_124_887_n1, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n5610, n579, n581, n590, n600,
         n6100, n620, n6300, n6500, n6600, n6700, n6800, n6900, n7000, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n17000, n17100,
         n17200, n17300, n17400, n17500, n17600, n17700, n17800, n17900,
         n18000, n18100, n18200, n18300, n18400, n18500, n18600, n18700,
         n18800, n18900, n19000, n19100, n19200, n19300, n19400, n19500,
         n19600, n19700, n19800, n19900, n20000, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n291, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n385, n387,
         n405, n406, n602, n603, n604, n605, n606, n607, n608, n609, n6101,
         n611, n612, n622, n623, n624, n625, n626, n627, n628, n629, n6301,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n6401, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n6501, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n6601, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n6701, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n6801, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n6901, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n7001, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n7101, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n7201, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n7301, n731, n732, n733, n734, n735, n736, n737, n738, n739, n7401,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n7501, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n7601, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n7701, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n7801, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n7901, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n8001, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n8101, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n8201, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n8301, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n8401, n841, n842, n843, n844, n845, n846, n847, n848, n849, n8501,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n8601, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n8801, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n8901, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n17001, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n17101, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n17201, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n17301, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n17401, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n17501, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n17601, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n17701, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n17801, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n17901, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n18001, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n18101, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n18201, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n18301, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n18401, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n18501, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n18601, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n18701, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n18801, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n18901, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n19001, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n19101, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n19201, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n19301, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n19401, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n19501, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n19601, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n19701, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n19801, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n19901, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n20001, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994;
  wire   [32:0] mul_operand_a_q;
  wire   [32:0] mul_operand_b_q;
  wire   [57:0] mult_result_w;
  wire   [31:1] q_mask_q;
  wire   [31:0] dividend_q;
  wire   [62:0] divisor_q;
  wire   [31:0] quotient_q;

  DFF_X1 mulhi_sel_q_reg ( .D(N89), .CK(clk_i), .Q(mulhi_sel_q), .QN(n2526) );
  SDFF_X1 mul_operand_a_q_reg_5_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[5]), 
        .CK(clk_i), .Q(mul_operand_a_q[5]), .QN(n1026) );
  DFF_X1 mul_operand_b_q_reg_2_ ( .D(N58), .CK(clk_i), .Q(mul_operand_b_q[2]), 
        .QN(n1008) );
  DFF_X1 mul_operand_b_q_reg_0_ ( .D(N56), .CK(clk_i), .Q(mul_operand_b_q[0]), 
        .QN(n1017) );
  DFF_X1 mul_busy_q_reg ( .D(n2499), .CK(clk_i), .Q(n2470), .QN(mul_busy_q) );
  DFF_X1 div_busy_q_reg ( .D(n578), .CK(clk_i), .Q(div_busy_q), .QN(n2473) );
  DFF_X1 invert_res_q_reg ( .D(n577), .CK(clk_i), .QN(n104) );
  DFF_X1 q_mask_q_reg_31_ ( .D(n576), .CK(clk_i), .Q(q_mask_q[31]), .QN(n2511)
         );
  DFF_X1 q_mask_q_reg_30_ ( .D(n545), .CK(clk_i), .Q(q_mask_q[30]), .QN(n2461)
         );
  DFF_X1 q_mask_q_reg_29_ ( .D(n546), .CK(clk_i), .Q(q_mask_q[29]), .QN(n2515)
         );
  DFF_X1 q_mask_q_reg_28_ ( .D(n547), .CK(clk_i), .Q(q_mask_q[28]), .QN(n2463)
         );
  DFF_X1 q_mask_q_reg_27_ ( .D(n548), .CK(clk_i), .Q(q_mask_q[27]), .QN(n2444)
         );
  DFF_X1 q_mask_q_reg_26_ ( .D(n549), .CK(clk_i), .Q(q_mask_q[26]), .QN(n2522)
         );
  DFF_X1 q_mask_q_reg_25_ ( .D(n550), .CK(clk_i), .Q(q_mask_q[25]), .QN(n2468)
         );
  DFF_X1 q_mask_q_reg_24_ ( .D(n551), .CK(clk_i), .Q(q_mask_q[24]), .QN(n2513)
         );
  DFF_X1 q_mask_q_reg_23_ ( .D(n552), .CK(clk_i), .Q(q_mask_q[23]), .QN(n2460)
         );
  DFF_X1 q_mask_q_reg_22_ ( .D(n553), .CK(clk_i), .Q(q_mask_q[22]), .QN(n2516)
         );
  DFF_X1 q_mask_q_reg_21_ ( .D(n554), .CK(clk_i), .Q(q_mask_q[21]), .QN(n2467)
         );
  DFF_X1 q_mask_q_reg_20_ ( .D(n555), .CK(clk_i), .Q(q_mask_q[20]), .QN(n2445)
         );
  DFF_X1 q_mask_q_reg_19_ ( .D(n556), .CK(clk_i), .Q(q_mask_q[19]), .QN(n2521)
         );
  DFF_X1 q_mask_q_reg_18_ ( .D(n557), .CK(clk_i), .Q(q_mask_q[18]), .QN(n2466)
         );
  DFF_X1 q_mask_q_reg_17_ ( .D(n558), .CK(clk_i), .Q(q_mask_q[17]), .QN(n2512)
         );
  DFF_X1 q_mask_q_reg_16_ ( .D(n559), .CK(clk_i), .Q(q_mask_q[16]), .QN(n2459)
         );
  DFF_X1 q_mask_q_reg_15_ ( .D(n560), .CK(clk_i), .Q(q_mask_q[15]), .QN(n2443)
         );
  DFF_X1 q_mask_q_reg_14_ ( .D(n561), .CK(clk_i), .Q(q_mask_q[14]), .QN(n2517)
         );
  DFF_X1 q_mask_q_reg_13_ ( .D(n562), .CK(clk_i), .Q(q_mask_q[13]), .QN(n2469)
         );
  DFF_X1 q_mask_q_reg_12_ ( .D(n563), .CK(clk_i), .Q(q_mask_q[12]), .QN(n2514)
         );
  DFF_X1 q_mask_q_reg_11_ ( .D(n564), .CK(clk_i), .Q(q_mask_q[11]), .QN(n2462)
         );
  DFF_X1 q_mask_q_reg_10_ ( .D(n565), .CK(clk_i), .Q(q_mask_q[10]), .QN(n2442)
         );
  DFF_X1 q_mask_q_reg_9_ ( .D(n566), .CK(clk_i), .Q(q_mask_q[9]), .QN(n2520)
         );
  DFF_X1 q_mask_q_reg_8_ ( .D(n567), .CK(clk_i), .Q(q_mask_q[8]), .QN(n2465)
         );
  DFF_X1 q_mask_q_reg_7_ ( .D(n568), .CK(clk_i), .QN(n6400) );
  DFF_X1 q_mask_q_reg_6_ ( .D(n569), .CK(clk_i), .Q(q_mask_q[6]), .QN(n2518)
         );
  DFF_X1 q_mask_q_reg_5_ ( .D(n570), .CK(clk_i), .Q(q_mask_q[5]), .QN(n2458)
         );
  DFF_X1 q_mask_q_reg_4_ ( .D(n571), .CK(clk_i), .Q(q_mask_q[4]), .QN(n2519)
         );
  DFF_X1 q_mask_q_reg_3_ ( .D(n572), .CK(clk_i), .Q(q_mask_q[3]), .QN(n2464)
         );
  DFF_X1 q_mask_q_reg_2_ ( .D(n573), .CK(clk_i), .Q(q_mask_q[2]), .QN(n2446)
         );
  DFF_X1 q_mask_q_reg_1_ ( .D(n574), .CK(clk_i), .Q(q_mask_q[1]), .QN(n2523)
         );
  DFF_X1 q_mask_q_reg_0_ ( .D(n5750), .CK(clk_i), .QN(n7100) );
  DFF_X1 dividend_q_reg_30_ ( .D(n482), .CK(clk_i), .Q(dividend_q[30]), .QN(
        n2492) );
  DFF_X1 dividend_q_reg_29_ ( .D(n483), .CK(clk_i), .Q(dividend_q[29]), .QN(
        n2452) );
  DFF_X1 dividend_q_reg_28_ ( .D(n484), .CK(clk_i), .Q(dividend_q[28]), .QN(
        n2496) );
  DFF_X1 dividend_q_reg_27_ ( .D(n485), .CK(clk_i), .Q(dividend_q[27]), .QN(
        n2456) );
  DFF_X1 dividend_q_reg_26_ ( .D(n486), .CK(clk_i), .Q(dividend_q[26]), .QN(
        n2489) );
  DFF_X1 dividend_q_reg_25_ ( .D(n487), .CK(clk_i), .Q(dividend_q[25]), .QN(
        n2454) );
  DFF_X1 dividend_q_reg_24_ ( .D(n488), .CK(clk_i), .Q(dividend_q[24]), .QN(
        n2498) );
  DFF_X1 dividend_q_reg_23_ ( .D(n489), .CK(clk_i), .Q(dividend_q[23]), .QN(
        n2453) );
  DFF_X1 dividend_q_reg_22_ ( .D(n490), .CK(clk_i), .Q(dividend_q[22]), .QN(
        n2490) );
  DFF_X1 dividend_q_reg_21_ ( .D(n491), .CK(clk_i), .Q(dividend_q[21]), .QN(
        n2451) );
  DFF_X1 dividend_q_reg_20_ ( .D(n492), .CK(clk_i), .Q(dividend_q[20]), .QN(
        n2497) );
  DFF_X1 dividend_q_reg_19_ ( .D(n493), .CK(clk_i), .Q(dividend_q[19]), .QN(
        n2457) );
  DFF_X1 dividend_q_reg_18_ ( .D(n494), .CK(clk_i), .Q(dividend_q[18]), .QN(
        n2491) );
  DFF_X1 dividend_q_reg_17_ ( .D(n495), .CK(clk_i), .Q(dividend_q[17]), .QN(
        n2455) );
  DFF_X1 dividend_q_reg_16_ ( .D(n496), .CK(clk_i), .Q(dividend_q[16]), .QN(
        n2493) );
  DFF_X1 dividend_q_reg_15_ ( .D(n497), .CK(clk_i), .Q(dividend_q[15]), .QN(
        n2475) );
  DFF_X1 dividend_q_reg_14_ ( .D(n498), .CK(clk_i), .Q(dividend_q[14]), .QN(
        n2480) );
  DFF_X1 dividend_q_reg_13_ ( .D(n499), .CK(clk_i), .Q(dividend_q[13]), .QN(
        n2449) );
  DFF_X1 dividend_q_reg_12_ ( .D(n500), .CK(clk_i), .Q(dividend_q[12]), .QN(
        n2477) );
  DFF_X1 dividend_q_reg_11_ ( .D(n501), .CK(clk_i), .Q(dividend_q[11]), .QN(
        n2479) );
  DFF_X1 dividend_q_reg_10_ ( .D(n502), .CK(clk_i), .Q(dividend_q[10]), .QN(
        n2476) );
  DFF_X1 dividend_q_reg_9_ ( .D(n503), .CK(clk_i), .Q(dividend_q[9]), .QN(
        n2450) );
  DFF_X1 dividend_q_reg_8_ ( .D(n504), .CK(clk_i), .Q(dividend_q[8]), .QN(
        n2478) );
  DFF_X1 dividend_q_reg_7_ ( .D(n505), .CK(clk_i), .Q(dividend_q[7]), .QN(
        n2484) );
  DFF_X1 dividend_q_reg_6_ ( .D(n506), .CK(clk_i), .Q(dividend_q[6]), .QN(
        n2482) );
  DFF_X1 dividend_q_reg_5_ ( .D(n507), .CK(clk_i), .Q(dividend_q[5]), .QN(
        n2485) );
  DFF_X1 dividend_q_reg_4_ ( .D(n508), .CK(clk_i), .Q(dividend_q[4]), .QN(
        n2481) );
  DFF_X1 dividend_q_reg_3_ ( .D(n509), .CK(clk_i), .Q(dividend_q[3]), .QN(
        n2471) );
  DFF_X1 dividend_q_reg_2_ ( .D(n510), .CK(clk_i), .Q(dividend_q[2]), .QN(
        n2447) );
  DFF_X1 dividend_q_reg_1_ ( .D(n511), .CK(clk_i), .Q(dividend_q[1]), .QN(
        n2448) );
  DFF_X1 dividend_q_reg_0_ ( .D(n512), .CK(clk_i), .Q(dividend_q[0]), .QN(
        n2472) );
  DFF_X1 dividend_q_reg_31_ ( .D(n513), .CK(clk_i), .Q(dividend_q[31]), .QN(
        n2524) );
  DFF_X1 quotient_q_reg_0_ ( .D(n480), .CK(clk_i), .Q(quotient_q[0]), .QN(n103) );
  DFF_X1 quotient_q_reg_1_ ( .D(n479), .CK(clk_i), .Q(quotient_q[1]), .QN(n102) );
  DFF_X1 quotient_q_reg_2_ ( .D(n478), .CK(clk_i), .Q(quotient_q[2]), .QN(n101) );
  DFF_X1 quotient_q_reg_3_ ( .D(n477), .CK(clk_i), .Q(quotient_q[3]), .QN(n100) );
  DFF_X1 quotient_q_reg_4_ ( .D(n476), .CK(clk_i), .Q(quotient_q[4]), .QN(n99)
         );
  DFF_X1 quotient_q_reg_5_ ( .D(n475), .CK(clk_i), .Q(quotient_q[5]), .QN(n98)
         );
  DFF_X1 quotient_q_reg_6_ ( .D(n474), .CK(clk_i), .Q(quotient_q[6]), .QN(n97)
         );
  DFF_X1 quotient_q_reg_7_ ( .D(n473), .CK(clk_i), .Q(quotient_q[7]), .QN(n96)
         );
  DFF_X1 quotient_q_reg_8_ ( .D(n472), .CK(clk_i), .Q(quotient_q[8]), .QN(n95)
         );
  DFF_X1 quotient_q_reg_9_ ( .D(n471), .CK(clk_i), .Q(quotient_q[9]), .QN(n94)
         );
  DFF_X1 quotient_q_reg_10_ ( .D(n470), .CK(clk_i), .Q(quotient_q[10]), .QN(
        n93) );
  DFF_X1 quotient_q_reg_11_ ( .D(n469), .CK(clk_i), .Q(quotient_q[11]), .QN(
        n92) );
  DFF_X1 quotient_q_reg_12_ ( .D(n468), .CK(clk_i), .Q(quotient_q[12]), .QN(
        n91) );
  DFF_X1 quotient_q_reg_13_ ( .D(n467), .CK(clk_i), .Q(quotient_q[13]), .QN(
        n90) );
  DFF_X1 quotient_q_reg_14_ ( .D(n466), .CK(clk_i), .Q(quotient_q[14]), .QN(
        n8900) );
  DFF_X1 quotient_q_reg_15_ ( .D(n465), .CK(clk_i), .Q(quotient_q[15]), .QN(
        n8800) );
  DFF_X1 quotient_q_reg_16_ ( .D(n464), .CK(clk_i), .Q(quotient_q[16]), .QN(
        n87) );
  DFF_X1 quotient_q_reg_17_ ( .D(n463), .CK(clk_i), .Q(quotient_q[17]), .QN(
        n8600) );
  DFF_X1 quotient_q_reg_18_ ( .D(n462), .CK(clk_i), .Q(quotient_q[18]), .QN(
        n8500) );
  DFF_X1 quotient_q_reg_19_ ( .D(n461), .CK(clk_i), .Q(quotient_q[19]), .QN(
        n8400) );
  DFF_X1 quotient_q_reg_20_ ( .D(n460), .CK(clk_i), .Q(quotient_q[20]), .QN(
        n8300) );
  DFF_X1 quotient_q_reg_21_ ( .D(n459), .CK(clk_i), .Q(quotient_q[21]), .QN(
        n8200) );
  DFF_X1 quotient_q_reg_22_ ( .D(n458), .CK(clk_i), .Q(quotient_q[22]), .QN(
        n8100) );
  DFF_X1 quotient_q_reg_23_ ( .D(n457), .CK(clk_i), .Q(quotient_q[23]), .QN(
        n8000) );
  DFF_X1 quotient_q_reg_24_ ( .D(n456), .CK(clk_i), .Q(quotient_q[24]), .QN(
        n7900) );
  DFF_X1 quotient_q_reg_25_ ( .D(n455), .CK(clk_i), .Q(quotient_q[25]), .QN(
        n7800) );
  DFF_X1 quotient_q_reg_26_ ( .D(n454), .CK(clk_i), .Q(quotient_q[26]), .QN(
        n7700) );
  DFF_X1 quotient_q_reg_27_ ( .D(n453), .CK(clk_i), .Q(quotient_q[27]), .QN(
        n7600) );
  DFF_X1 quotient_q_reg_28_ ( .D(n452), .CK(clk_i), .Q(quotient_q[28]), .QN(
        n7500) );
  DFF_X1 quotient_q_reg_29_ ( .D(n451), .CK(clk_i), .Q(quotient_q[29]), .QN(
        n7400) );
  DFF_X1 quotient_q_reg_30_ ( .D(n450), .CK(clk_i), .Q(quotient_q[30]), .QN(
        n7300) );
  DFF_X1 quotient_q_reg_31_ ( .D(n481), .CK(clk_i), .Q(quotient_q[31]), .QN(
        n7200) );
  DFF_X1 divisor_q_reg_62_ ( .D(n386), .CK(clk_i), .QN(divisor_q[62]) );
  DFF_X1 divisor_q_reg_30_ ( .D(n290), .CK(clk_i), .QN(divisor_q[30]) );
  DFF_X1 divisor_q_reg_29_ ( .D(n292), .CK(clk_i), .QN(divisor_q[29]) );
  DFF_X1 divisor_q_reg_28_ ( .D(n293), .CK(clk_i), .Q(n2506), .QN(
        divisor_q[28]) );
  DFF_X1 divisor_q_reg_27_ ( .D(n294), .CK(clk_i), .Q(n2502), .QN(
        divisor_q[27]) );
  DFF_X1 divisor_q_reg_26_ ( .D(n295), .CK(clk_i), .QN(divisor_q[26]) );
  DFF_X1 divisor_q_reg_25_ ( .D(n296), .CK(clk_i), .QN(divisor_q[25]) );
  DFF_X1 divisor_q_reg_24_ ( .D(n297), .CK(clk_i), .Q(n2507), .QN(
        divisor_q[24]) );
  DFF_X1 divisor_q_reg_23_ ( .D(n298), .CK(clk_i), .QN(divisor_q[23]) );
  DFF_X1 divisor_q_reg_22_ ( .D(n299), .CK(clk_i), .QN(divisor_q[22]) );
  DFF_X1 divisor_q_reg_21_ ( .D(n300), .CK(clk_i), .QN(divisor_q[21]) );
  DFF_X1 divisor_q_reg_20_ ( .D(n301), .CK(clk_i), .Q(n2505), .QN(
        divisor_q[20]) );
  DFF_X1 divisor_q_reg_19_ ( .D(n302), .CK(clk_i), .Q(n2501), .QN(
        divisor_q[19]) );
  DFF_X1 divisor_q_reg_18_ ( .D(n303), .CK(clk_i), .QN(divisor_q[18]) );
  DFF_X1 divisor_q_reg_17_ ( .D(n304), .CK(clk_i), .QN(divisor_q[17]) );
  DFF_X1 divisor_q_reg_16_ ( .D(n305), .CK(clk_i), .QN(divisor_q[16]) );
  DFF_X1 divisor_q_reg_15_ ( .D(n306), .CK(clk_i), .Q(n2488), .QN(
        divisor_q[15]) );
  DFF_X1 divisor_q_reg_14_ ( .D(n307), .CK(clk_i), .Q(n2509), .QN(
        divisor_q[14]) );
  DFF_X1 divisor_q_reg_13_ ( .D(n308), .CK(clk_i), .QN(divisor_q[13]) );
  DFF_X1 divisor_q_reg_12_ ( .D(n309), .CK(clk_i), .QN(divisor_q[12]) );
  DFF_X1 divisor_q_reg_11_ ( .D(n310), .CK(clk_i), .Q(n2508), .QN(
        divisor_q[11]) );
  DFF_X1 divisor_q_reg_10_ ( .D(n311), .CK(clk_i), .QN(divisor_q[10]) );
  DFF_X1 divisor_q_reg_9_ ( .D(n312), .CK(clk_i), .QN(divisor_q[9]) );
  DFF_X1 divisor_q_reg_8_ ( .D(n313), .CK(clk_i), .Q(n2504), .QN(divisor_q[8])
         );
  DFF_X1 divisor_q_reg_7_ ( .D(n314), .CK(clk_i), .Q(n2495), .QN(divisor_q[7])
         );
  DFF_X1 divisor_q_reg_6_ ( .D(n315), .CK(clk_i), .QN(divisor_q[6]) );
  DFF_X1 divisor_q_reg_5_ ( .D(n316), .CK(clk_i), .Q(n2494), .QN(divisor_q[5])
         );
  DFF_X1 divisor_q_reg_4_ ( .D(n317), .CK(clk_i), .QN(divisor_q[4]) );
  DFF_X1 divisor_q_reg_3_ ( .D(n318), .CK(clk_i), .Q(n2503), .QN(divisor_q[3])
         );
  DFF_X1 divisor_q_reg_2_ ( .D(n319), .CK(clk_i), .QN(divisor_q[2]) );
  DFF_X1 divisor_q_reg_1_ ( .D(n320), .CK(clk_i), .Q(n2510), .QN(divisor_q[1])
         );
  DFF_X1 divisor_q_reg_0_ ( .D(n321), .CK(clk_i), .Q(n2474), .QN(divisor_q[0])
         );
  DFF_X1 div_inst_q_reg ( .D(n449), .CK(clk_i), .Q(div_inst_q), .QN(n2483) );
  DFF_X1 result_q_reg_29_ ( .D(n446), .CK(clk_i), .Q(result_o[29]) );
  DFF_X1 result_q_reg_2_ ( .D(n419), .CK(clk_i), .Q(result_o[2]), .QN(n2527)
         );
  DFF_X1 result_q_reg_1_ ( .D(n418), .CK(clk_i), .Q(result_o[1]), .QN(n2525)
         );
  HA_X1 sub_x_9_U31 ( .A(n2535), .B(n2536), .CO(sub_x_9_n30), .S(N170) );
  HA_X1 sub_x_9_U30 ( .A(sub_x_9_n30), .B(n2537), .CO(sub_x_9_n29), .S(N171)
         );
  HA_X1 sub_x_9_U29 ( .A(sub_x_9_n29), .B(n2538), .CO(sub_x_9_n28), .S(N172)
         );
  HA_X1 sub_x_9_U28 ( .A(sub_x_9_n28), .B(n2539), .CO(sub_x_9_n27), .S(N173)
         );
  HA_X1 sub_x_9_U27 ( .A(sub_x_9_n27), .B(n2540), .CO(sub_x_9_n26), .S(N174)
         );
  HA_X1 sub_x_9_U26 ( .A(sub_x_9_n26), .B(n2541), .CO(sub_x_9_n25), .S(N175)
         );
  HA_X1 sub_x_9_U25 ( .A(sub_x_9_n25), .B(n2542), .CO(sub_x_9_n24), .S(N176)
         );
  HA_X1 sub_x_9_U24 ( .A(sub_x_9_n24), .B(n2543), .CO(sub_x_9_n23), .S(N177)
         );
  HA_X1 sub_x_9_U23 ( .A(sub_x_9_n23), .B(n2544), .CO(sub_x_9_n22), .S(N178)
         );
  HA_X1 sub_x_9_U22 ( .A(sub_x_9_n22), .B(n2545), .CO(sub_x_9_n21), .S(N179)
         );
  HA_X1 sub_x_9_U21 ( .A(sub_x_9_n21), .B(n2546), .CO(sub_x_9_n20), .S(N180)
         );
  HA_X1 sub_x_9_U20 ( .A(sub_x_9_n20), .B(n2547), .CO(sub_x_9_n19), .S(N181)
         );
  HA_X1 sub_x_9_U19 ( .A(sub_x_9_n19), .B(n2548), .CO(sub_x_9_n18), .S(N182)
         );
  HA_X1 sub_x_9_U18 ( .A(sub_x_9_n18), .B(n2549), .CO(sub_x_9_n17), .S(N183)
         );
  HA_X1 sub_x_9_U17 ( .A(sub_x_9_n17), .B(n2550), .CO(sub_x_9_n16), .S(N184)
         );
  HA_X1 sub_x_9_U16 ( .A(sub_x_9_n16), .B(n2551), .CO(sub_x_9_n15), .S(N185)
         );
  HA_X1 sub_x_9_U15 ( .A(sub_x_9_n15), .B(n2552), .CO(sub_x_9_n14), .S(N186)
         );
  HA_X1 sub_x_9_U14 ( .A(sub_x_9_n14), .B(n2553), .CO(sub_x_9_n13), .S(N187)
         );
  HA_X1 sub_x_9_U13 ( .A(sub_x_9_n13), .B(n2554), .CO(sub_x_9_n12), .S(N188)
         );
  HA_X1 sub_x_9_U12 ( .A(sub_x_9_n12), .B(n2555), .CO(sub_x_9_n11), .S(N189)
         );
  HA_X1 sub_x_9_U11 ( .A(sub_x_9_n11), .B(n2556), .CO(sub_x_9_n10), .S(N190)
         );
  HA_X1 sub_x_9_U10 ( .A(sub_x_9_n10), .B(n2557), .CO(sub_x_9_n9), .S(N191) );
  HA_X1 sub_x_9_U9 ( .A(sub_x_9_n9), .B(n2558), .CO(sub_x_9_n8), .S(N192) );
  HA_X1 sub_x_9_U8 ( .A(sub_x_9_n8), .B(n2559), .CO(sub_x_9_n7), .S(N193) );
  HA_X1 sub_x_9_U7 ( .A(sub_x_9_n7), .B(n2560), .CO(sub_x_9_n6), .S(N194) );
  HA_X1 sub_x_9_U6 ( .A(sub_x_9_n6), .B(n2561), .CO(sub_x_9_n5), .S(N195) );
  HA_X1 sub_x_9_U5 ( .A(sub_x_9_n5), .B(n2562), .CO(sub_x_9_n4), .S(N196) );
  HA_X1 sub_x_9_U4 ( .A(sub_x_9_n4), .B(n2563), .CO(sub_x_9_n3), .S(N197) );
  HA_X1 sub_x_9_U3 ( .A(sub_x_9_n3), .B(n2564), .CO(sub_x_9_n2), .S(N198) );
  HA_X1 sub_x_9_U2 ( .A(sub_x_9_n2), .B(n2565), .CO(sub_x_9_n1), .S(N199) );
  HA_X1 DP_OP_63J3_127_9516_U31 ( .A(n2746), .B(n2743), .CO(
        DP_OP_63J3_127_9516_n30), .S(C22_DATA3_1) );
  HA_X1 DP_OP_63J3_127_9516_U30 ( .A(DP_OP_63J3_127_9516_n30), .B(n2740), .CO(
        DP_OP_63J3_127_9516_n29), .S(C22_DATA3_2) );
  HA_X1 DP_OP_63J3_127_9516_U29 ( .A(DP_OP_63J3_127_9516_n29), .B(n2739), .CO(
        DP_OP_63J3_127_9516_n28), .S(C22_DATA3_3) );
  HA_X1 DP_OP_63J3_127_9516_U28 ( .A(DP_OP_63J3_127_9516_n28), .B(n2738), .CO(
        DP_OP_63J3_127_9516_n27), .S(C22_DATA3_4) );
  HA_X1 DP_OP_63J3_127_9516_U27 ( .A(DP_OP_63J3_127_9516_n27), .B(n2737), .CO(
        DP_OP_63J3_127_9516_n26), .S(C22_DATA3_5) );
  HA_X1 DP_OP_63J3_127_9516_U26 ( .A(DP_OP_63J3_127_9516_n26), .B(n2736), .CO(
        DP_OP_63J3_127_9516_n25), .S(C22_DATA3_6) );
  HA_X1 DP_OP_63J3_127_9516_U25 ( .A(DP_OP_63J3_127_9516_n25), .B(n2735), .CO(
        DP_OP_63J3_127_9516_n24), .S(C22_DATA3_7) );
  HA_X1 DP_OP_63J3_127_9516_U24 ( .A(DP_OP_63J3_127_9516_n24), .B(n2734), .CO(
        DP_OP_63J3_127_9516_n23), .S(C22_DATA3_8) );
  HA_X1 DP_OP_63J3_127_9516_U23 ( .A(DP_OP_63J3_127_9516_n23), .B(n2733), .CO(
        DP_OP_63J3_127_9516_n22), .S(C22_DATA3_9) );
  HA_X1 DP_OP_63J3_127_9516_U22 ( .A(DP_OP_63J3_127_9516_n22), .B(n2732), .CO(
        DP_OP_63J3_127_9516_n21), .S(C22_DATA3_10) );
  HA_X1 DP_OP_63J3_127_9516_U21 ( .A(DP_OP_63J3_127_9516_n21), .B(n2731), .CO(
        DP_OP_63J3_127_9516_n20), .S(C22_DATA3_11) );
  HA_X1 DP_OP_63J3_127_9516_U20 ( .A(DP_OP_63J3_127_9516_n20), .B(n2730), .CO(
        DP_OP_63J3_127_9516_n19), .S(C22_DATA3_12) );
  HA_X1 DP_OP_63J3_127_9516_U19 ( .A(DP_OP_63J3_127_9516_n19), .B(n2729), .CO(
        DP_OP_63J3_127_9516_n18), .S(C22_DATA3_13) );
  HA_X1 DP_OP_63J3_127_9516_U18 ( .A(DP_OP_63J3_127_9516_n18), .B(n2728), .CO(
        DP_OP_63J3_127_9516_n17), .S(C22_DATA3_14) );
  HA_X1 DP_OP_63J3_127_9516_U17 ( .A(DP_OP_63J3_127_9516_n17), .B(n2727), .CO(
        DP_OP_63J3_127_9516_n16), .S(C22_DATA3_15) );
  HA_X1 DP_OP_63J3_127_9516_U16 ( .A(DP_OP_63J3_127_9516_n16), .B(n2726), .CO(
        DP_OP_63J3_127_9516_n15), .S(C22_DATA3_16) );
  HA_X1 DP_OP_63J3_127_9516_U15 ( .A(DP_OP_63J3_127_9516_n15), .B(n2725), .CO(
        DP_OP_63J3_127_9516_n14), .S(C22_DATA3_17) );
  HA_X1 DP_OP_63J3_127_9516_U14 ( .A(DP_OP_63J3_127_9516_n14), .B(n2724), .CO(
        DP_OP_63J3_127_9516_n13), .S(C22_DATA3_18) );
  HA_X1 DP_OP_63J3_127_9516_U13 ( .A(DP_OP_63J3_127_9516_n13), .B(n2723), .CO(
        DP_OP_63J3_127_9516_n12), .S(C22_DATA3_19) );
  HA_X1 DP_OP_63J3_127_9516_U12 ( .A(DP_OP_63J3_127_9516_n12), .B(n2722), .CO(
        DP_OP_63J3_127_9516_n11), .S(C22_DATA3_20) );
  HA_X1 DP_OP_63J3_127_9516_U11 ( .A(DP_OP_63J3_127_9516_n11), .B(n2721), .CO(
        DP_OP_63J3_127_9516_n10), .S(C22_DATA3_21) );
  HA_X1 DP_OP_63J3_127_9516_U10 ( .A(DP_OP_63J3_127_9516_n10), .B(n2720), .CO(
        DP_OP_63J3_127_9516_n9), .S(C22_DATA3_22) );
  HA_X1 DP_OP_63J3_127_9516_U9 ( .A(DP_OP_63J3_127_9516_n9), .B(n2719), .CO(
        DP_OP_63J3_127_9516_n8), .S(C22_DATA3_23) );
  HA_X1 DP_OP_63J3_127_9516_U8 ( .A(DP_OP_63J3_127_9516_n8), .B(n2718), .CO(
        DP_OP_63J3_127_9516_n7), .S(C22_DATA3_24) );
  HA_X1 DP_OP_63J3_127_9516_U7 ( .A(DP_OP_63J3_127_9516_n7), .B(n2717), .CO(
        DP_OP_63J3_127_9516_n6), .S(C22_DATA3_25) );
  HA_X1 DP_OP_63J3_127_9516_U6 ( .A(DP_OP_63J3_127_9516_n6), .B(n2716), .CO(
        DP_OP_63J3_127_9516_n5), .S(C22_DATA3_26) );
  HA_X1 DP_OP_63J3_127_9516_U5 ( .A(DP_OP_63J3_127_9516_n5), .B(n2715), .CO(
        DP_OP_63J3_127_9516_n4), .S(C22_DATA3_27) );
  HA_X1 DP_OP_63J3_127_9516_U4 ( .A(DP_OP_63J3_127_9516_n4), .B(n2714), .CO(
        DP_OP_63J3_127_9516_n3), .S(C22_DATA3_28) );
  HA_X1 DP_OP_63J3_127_9516_U3 ( .A(DP_OP_63J3_127_9516_n3), .B(n2713), .CO(
        DP_OP_63J3_127_9516_n2), .S(C22_DATA3_29) );
  HA_X1 DP_OP_63J3_127_9516_U2 ( .A(DP_OP_63J3_127_9516_n2), .B(n2712), .CO(
        DP_OP_63J3_127_9516_n1), .S(C22_DATA3_30) );
  DFF_X1 mul_operand_a_q_reg_1_ ( .D(n2530), .CK(clk_i), .Q(mul_operand_a_q[1]), .QN(n1014) );
  FA_X1 mult_x_6_U2045 ( .A(n1015), .B(mul_operand_b_q[2]), .CI(mult_x_6_n1070), .CO(mult_x_6_n1069), .S(mult_x_6_n1102) );
  FA_X1 mult_x_6_U2026 ( .A(mul_operand_b_q[20]), .B(mul_operand_b_q[21]), 
        .CI(mult_x_6_n1051), .CO(mult_x_6_n1050), .S(mult_x_6_n1083) );
  FA_X1 mult_x_6_U2025 ( .A(mul_operand_b_q[21]), .B(mul_operand_b_q[22]), 
        .CI(mult_x_6_n1050), .CO(mult_x_6_n1049), .S(mult_x_6_n1082) );
  FA_X1 mult_x_6_U2022 ( .A(n2183), .B(mul_operand_b_q[25]), .CI(
        mult_x_6_n1047), .CO(mult_x_6_n1046), .S(mult_x_6_n1079) );
  FA_X1 mult_x_6_U2015 ( .A(n2179), .B(n2177), .CI(mult_x_6_n1040), .CO(
        mult_x_6_n1071), .S(mult_x_6_n1072) );
  HA_X1 mult_x_6_U669 ( .A(mult_x_6_n1413), .B(n2174), .CO(mult_x_6_n988), .S(
        mult_x_6_n989) );
  FA_X1 mult_x_6_U666 ( .A(mult_x_6_n1444), .B(mult_x_6_n985), .CI(
        mult_x_6_n986), .CO(mult_x_6_n982), .S(mult_x_6_n983) );
  FA_X1 mult_x_6_U662 ( .A(mult_x_6_n1410), .B(mult_x_6_n977), .CI(
        mult_x_6_n980), .CO(mult_x_6_n974), .S(mult_x_6_n975) );
  FA_X1 mult_x_6_U661 ( .A(mult_x_6_n1442), .B(mult_x_6_n975), .CI(
        mult_x_6_n978), .CO(mult_x_6_n972), .S(mult_x_6_n973) );
  HA_X1 mult_x_6_U657 ( .A(mult_x_6_n970), .B(mult_x_6_n1376), .CO(
        mult_x_6_n964), .S(mult_x_6_n965) );
  FA_X1 mult_x_6_U653 ( .A(mult_x_6_n1375), .B(mult_x_6_n959), .CI(
        mult_x_6_n964), .CO(mult_x_6_n956), .S(mult_x_6_n957) );
  FA_X1 mult_x_6_U652 ( .A(mult_x_6_n1407), .B(mult_x_6_n957), .CI(
        mult_x_6_n962), .CO(mult_x_6_n954), .S(mult_x_6_n955) );
  HA_X1 mult_x_6_U646 ( .A(mult_x_6_n950), .B(mult_x_6_n1341), .CO(
        mult_x_6_n942), .S(mult_x_6_n943) );
  FA_X1 mult_x_6_U641 ( .A(mult_x_6_n1340), .B(mult_x_6_n935), .CI(
        mult_x_6_n942), .CO(mult_x_6_n932), .S(mult_x_6_n933) );
  FA_X1 mult_x_6_U640 ( .A(mult_x_6_n1372), .B(mult_x_6_n933), .CI(
        mult_x_6_n940), .CO(mult_x_6_n930), .S(mult_x_6_n931) );
  FA_X1 mult_x_6_U639 ( .A(mult_x_6_n1404), .B(mult_x_6_n931), .CI(
        mult_x_6_n938), .CO(mult_x_6_n928), .S(mult_x_6_n929) );
  FA_X1 mult_x_6_U636 ( .A(mult_x_6_n1339), .B(mult_x_6_n925), .CI(
        mult_x_6_n932), .CO(mult_x_6_n922), .S(mult_x_6_n923) );
  FA_X1 mult_x_6_U635 ( .A(mult_x_6_n1371), .B(mult_x_6_n923), .CI(
        mult_x_6_n930), .CO(mult_x_6_n920), .S(mult_x_6_n921) );
  HA_X1 mult_x_6_U632 ( .A(mult_x_6_n924), .B(mult_x_6_n1306), .CO(
        mult_x_6_n914), .S(mult_x_6_n915) );
  FA_X1 mult_x_6_U631 ( .A(mult_x_6_n1338), .B(mult_x_6_n915), .CI(
        mult_x_6_n922), .CO(mult_x_6_n912), .S(mult_x_6_n913) );
  HA_X1 mult_x_6_U627 ( .A(mult_x_6_n1273), .B(n2170), .CO(mult_x_6_n904), .S(
        mult_x_6_n905) );
  FA_X1 mult_x_6_U626 ( .A(mult_x_6_n1305), .B(mult_x_6_n905), .CI(
        mult_x_6_n914), .CO(mult_x_6_n902), .S(mult_x_6_n903) );
  FA_X1 mult_x_6_U625 ( .A(mult_x_6_n1337), .B(mult_x_6_n903), .CI(
        mult_x_6_n912), .CO(mult_x_6_n900), .S(mult_x_6_n901) );
  FA_X1 mult_x_6_U623 ( .A(mult_x_6_n1401), .B(mult_x_6_n899), .CI(
        mult_x_6_n908), .CO(mult_x_6_n896), .S(mult_x_6_n897) );
  FA_X1 mult_x_6_U622 ( .A(mult_x_6_n1433), .B(mult_x_6_n897), .CI(
        mult_x_6_n906), .CO(mult_x_6_n894), .S(mult_x_6_n895) );
  HA_X1 mult_x_6_U621 ( .A(mult_x_6_n904), .B(mult_x_6_n1272), .CO(
        mult_x_6_n892), .S(mult_x_6_n893) );
  FA_X1 mult_x_6_U620 ( .A(mult_x_6_n1304), .B(mult_x_6_n893), .CI(
        mult_x_6_n902), .CO(mult_x_6_n890), .S(mult_x_6_n891) );
  FA_X1 mult_x_6_U619 ( .A(mult_x_6_n1336), .B(mult_x_6_n891), .CI(
        mult_x_6_n900), .CO(mult_x_6_n888), .S(mult_x_6_n889) );
  FA_X1 mult_x_6_U617 ( .A(mult_x_6_n1400), .B(mult_x_6_n887), .CI(
        mult_x_6_n896), .CO(mult_x_6_n884), .S(mult_x_6_n885) );
  FA_X1 mult_x_6_U616 ( .A(mult_x_6_n1432), .B(mult_x_6_n885), .CI(
        mult_x_6_n894), .CO(mult_x_6_n882), .S(mult_x_6_n883) );
  HA_X1 mult_x_6_U615 ( .A(mult_x_6_n892), .B(mult_x_6_n1271), .CO(
        mult_x_6_n880), .S(mult_x_6_n881) );
  FA_X1 mult_x_6_U614 ( .A(mult_x_6_n1303), .B(mult_x_6_n881), .CI(
        mult_x_6_n890), .CO(mult_x_6_n878), .S(mult_x_6_n879) );
  FA_X1 mult_x_6_U613 ( .A(mult_x_6_n1335), .B(mult_x_6_n879), .CI(
        mult_x_6_n888), .CO(mult_x_6_n876), .S(mult_x_6_n877) );
  FA_X1 mult_x_6_U612 ( .A(mult_x_6_n1367), .B(mult_x_6_n877), .CI(
        mult_x_6_n886), .CO(mult_x_6_n874), .S(mult_x_6_n875) );
  HA_X1 mult_x_6_U609 ( .A(mult_x_6_n1238), .B(mul_operand_a_q[23]), .CO(
        mult_x_6_n868), .S(mult_x_6_n869) );
  FA_X1 mult_x_6_U608 ( .A(mult_x_6_n1270), .B(mult_x_6_n869), .CI(
        mult_x_6_n880), .CO(mult_x_6_n866), .S(mult_x_6_n867) );
  FA_X1 mult_x_6_U607 ( .A(mult_x_6_n1302), .B(mult_x_6_n867), .CI(
        mult_x_6_n878), .CO(mult_x_6_n864), .S(mult_x_6_n865) );
  FA_X1 mult_x_6_U606 ( .A(mult_x_6_n1334), .B(mult_x_6_n865), .CI(
        mult_x_6_n876), .CO(mult_x_6_n862), .S(mult_x_6_n863) );
  FA_X1 mult_x_6_U605 ( .A(mult_x_6_n1366), .B(mult_x_6_n863), .CI(
        mult_x_6_n874), .CO(mult_x_6_n860), .S(mult_x_6_n861) );
  HA_X1 mult_x_6_U602 ( .A(mult_x_6_n868), .B(mult_x_6_n1237), .CO(
        mult_x_6_n854), .S(mult_x_6_n855) );
  FA_X1 mult_x_6_U601 ( .A(mult_x_6_n1269), .B(mult_x_6_n855), .CI(
        mult_x_6_n866), .CO(mult_x_6_n852), .S(mult_x_6_n853) );
  FA_X1 mult_x_6_U600 ( .A(mult_x_6_n1301), .B(mult_x_6_n853), .CI(
        mult_x_6_n864), .CO(mult_x_6_n850), .S(mult_x_6_n851) );
  FA_X1 mult_x_6_U599 ( .A(mult_x_6_n1333), .B(mult_x_6_n851), .CI(
        mult_x_6_n862), .CO(mult_x_6_n848), .S(mult_x_6_n849) );
  HA_X1 mult_x_6_U595 ( .A(mult_x_6_n854), .B(mult_x_6_n1236), .CO(
        mult_x_6_n840), .S(mult_x_6_n841) );
  FA_X1 mult_x_6_U594 ( .A(mult_x_6_n1268), .B(mult_x_6_n841), .CI(
        mult_x_6_n852), .CO(mult_x_6_n838), .S(mult_x_6_n839) );
  FA_X1 mult_x_6_U593 ( .A(mult_x_6_n1300), .B(mult_x_6_n839), .CI(
        mult_x_6_n850), .CO(mult_x_6_n836), .S(mult_x_6_n837) );
  FA_X1 mult_x_6_U590 ( .A(mult_x_6_n1396), .B(mult_x_6_n833), .CI(
        mult_x_6_n844), .CO(mult_x_6_n830), .S(mult_x_6_n831) );
  FA_X1 mult_x_6_U589 ( .A(mult_x_6_n1428), .B(mult_x_6_n831), .CI(
        mult_x_6_n842), .CO(mult_x_6_n828), .S(mult_x_6_n829) );
  HA_X1 mult_x_6_U588 ( .A(mult_x_6_n1203), .B(mul_operand_a_q[26]), .CO(
        mult_x_6_n826), .S(mult_x_6_n827) );
  FA_X1 mult_x_6_U587 ( .A(mult_x_6_n1235), .B(mult_x_6_n827), .CI(
        mult_x_6_n840), .CO(mult_x_6_n824), .S(mult_x_6_n825) );
  FA_X1 mult_x_6_U586 ( .A(mult_x_6_n1267), .B(mult_x_6_n825), .CI(
        mult_x_6_n838), .CO(mult_x_6_n822), .S(mult_x_6_n823) );
  FA_X1 mult_x_6_U585 ( .A(mult_x_6_n1299), .B(mult_x_6_n823), .CI(
        mult_x_6_n836), .CO(mult_x_6_n820), .S(mult_x_6_n821) );
  HA_X1 mult_x_6_U580 ( .A(mult_x_6_n826), .B(mult_x_6_n1202), .CO(
        mult_x_6_n810), .S(mult_x_6_n811) );
  FA_X1 mult_x_6_U579 ( .A(mult_x_6_n1234), .B(mult_x_6_n811), .CI(
        mult_x_6_n824), .CO(mult_x_6_n808), .S(mult_x_6_n809) );
  FA_X1 mult_x_6_U578 ( .A(mult_x_6_n1266), .B(mult_x_6_n809), .CI(
        mult_x_6_n822), .CO(mult_x_6_n806), .S(mult_x_6_n807) );
  FA_X1 mult_x_6_U577 ( .A(mult_x_6_n1298), .B(mult_x_6_n807), .CI(
        mult_x_6_n820), .CO(mult_x_6_n804), .S(mult_x_6_n805) );
  HA_X1 mult_x_6_U572 ( .A(mult_x_6_n810), .B(mult_x_6_n1201), .CO(
        mult_x_6_n794), .S(mult_x_6_n795) );
  FA_X1 mult_x_6_U571 ( .A(mult_x_6_n1233), .B(mult_x_6_n795), .CI(
        mult_x_6_n808), .CO(mult_x_6_n792), .S(mult_x_6_n793) );
  FA_X1 mult_x_6_U570 ( .A(mult_x_6_n1265), .B(mult_x_6_n793), .CI(
        mult_x_6_n806), .CO(mult_x_6_n790), .S(mult_x_6_n791) );
  FA_X1 mult_x_6_U569 ( .A(mult_x_6_n1297), .B(mult_x_6_n791), .CI(
        mult_x_6_n804), .CO(mult_x_6_n788), .S(mult_x_6_n789) );
  HA_X1 mult_x_6_U564 ( .A(mult_x_6_n1168), .B(mul_operand_a_q[29]), .CO(
        mult_x_6_n778), .S(mult_x_6_n779) );
  FA_X1 mult_x_6_U563 ( .A(mult_x_6_n1200), .B(mult_x_6_n779), .CI(
        mult_x_6_n794), .CO(mult_x_6_n776), .S(mult_x_6_n777) );
  FA_X1 mult_x_6_U562 ( .A(mult_x_6_n1232), .B(mult_x_6_n777), .CI(
        mult_x_6_n792), .CO(mult_x_6_n774), .S(mult_x_6_n775) );
  FA_X1 mult_x_6_U561 ( .A(mult_x_6_n1264), .B(mult_x_6_n775), .CI(
        mult_x_6_n790), .CO(mult_x_6_n772), .S(mult_x_6_n773) );
  FA_X1 mult_x_6_U560 ( .A(mult_x_6_n1296), .B(mult_x_6_n773), .CI(
        mult_x_6_n788), .CO(mult_x_6_n770), .S(mult_x_6_n771) );
  FA_X1 mult_x_6_U558 ( .A(mult_x_6_n1360), .B(mult_x_6_n769), .CI(
        mult_x_6_n784), .CO(mult_x_6_n766), .S(mult_x_6_n767) );
  FA_X1 mult_x_6_U557 ( .A(mult_x_6_n1392), .B(mult_x_6_n767), .CI(
        mult_x_6_n782), .CO(mult_x_6_n764), .S(mult_x_6_n765) );
  HA_X1 mult_x_6_U555 ( .A(mult_x_6_n778), .B(mult_x_6_n1167), .CO(
        mult_x_6_n760), .S(mult_x_6_n761) );
  FA_X1 mult_x_6_U554 ( .A(mult_x_6_n1199), .B(mult_x_6_n761), .CI(
        mult_x_6_n776), .CO(mult_x_6_n758), .S(mult_x_6_n759) );
  FA_X1 mult_x_6_U553 ( .A(mult_x_6_n1231), .B(mult_x_6_n759), .CI(
        mult_x_6_n774), .CO(mult_x_6_n756), .S(mult_x_6_n757) );
  FA_X1 mult_x_6_U552 ( .A(mult_x_6_n1263), .B(mult_x_6_n757), .CI(
        mult_x_6_n772), .CO(mult_x_6_n754), .S(mult_x_6_n755) );
  FA_X1 mult_x_6_U551 ( .A(mult_x_6_n1295), .B(mult_x_6_n755), .CI(
        mult_x_6_n770), .CO(mult_x_6_n752), .S(mult_x_6_n753) );
  FA_X1 mult_x_6_U550 ( .A(mult_x_6_n1327), .B(mult_x_6_n753), .CI(
        mult_x_6_n768), .CO(mult_x_6_n750), .S(mult_x_6_n751) );
  FA_X1 mult_x_6_U548 ( .A(mult_x_6_n1391), .B(mult_x_6_n749), .CI(
        mult_x_6_n764), .CO(mult_x_6_n746), .S(mult_x_6_n747) );
  FA_X1 mult_x_6_U547 ( .A(mult_x_6_n1423), .B(mult_x_6_n747), .CI(
        mult_x_6_n762), .CO(mult_x_6_n744), .S(mult_x_6_n745) );
  HA_X1 mult_x_6_U546 ( .A(mult_x_6_n760), .B(mult_x_6_n1166), .CO(
        mult_x_6_n742), .S(mult_x_6_n743) );
  FA_X1 mult_x_6_U545 ( .A(mult_x_6_n1198), .B(mult_x_6_n743), .CI(
        mult_x_6_n758), .CO(mult_x_6_n740), .S(mult_x_6_n741) );
  FA_X1 mult_x_6_U544 ( .A(mult_x_6_n1230), .B(mult_x_6_n741), .CI(
        mult_x_6_n756), .CO(mult_x_6_n738), .S(mult_x_6_n739) );
  FA_X1 mult_x_6_U543 ( .A(mult_x_6_n1262), .B(mult_x_6_n739), .CI(
        mult_x_6_n754), .CO(mult_x_6_n736), .S(mult_x_6_n737) );
  HA_X1 mult_x_6_U537 ( .A(mult_x_6_n1133), .B(mul_operand_a_q[32]), .CO(
        mult_x_6_n724), .S(mult_x_6_n725) );
  FA_X1 mult_x_6_U536 ( .A(mult_x_6_n1165), .B(mult_x_6_n725), .CI(
        mult_x_6_n742), .CO(mult_x_6_n722), .S(mult_x_6_n723) );
  FA_X1 mult_x_6_U535 ( .A(mult_x_6_n1197), .B(mult_x_6_n723), .CI(
        mult_x_6_n740), .CO(mult_x_6_n720), .S(mult_x_6_n721) );
  FA_X1 mult_x_6_U534 ( .A(mult_x_6_n1229), .B(mult_x_6_n721), .CI(
        mult_x_6_n738), .CO(mult_x_6_n718), .S(mult_x_6_n719) );
  FA_X1 mult_x_6_U533 ( .A(mult_x_6_n1261), .B(mult_x_6_n719), .CI(
        mult_x_6_n736), .CO(mult_x_6_n716), .S(mult_x_6_n717) );
  FA_X1 mult_x_6_U532 ( .A(mult_x_6_n1293), .B(mult_x_6_n717), .CI(
        mult_x_6_n734), .CO(mult_x_6_n714), .S(mult_x_6_n715) );
  FA_X1 mult_x_6_U531 ( .A(mult_x_6_n1325), .B(mult_x_6_n715), .CI(
        mult_x_6_n732), .CO(mult_x_6_n712), .S(mult_x_6_n713) );
  FA_X1 mult_x_6_U530 ( .A(mult_x_6_n1357), .B(mult_x_6_n713), .CI(
        mult_x_6_n730), .CO(mult_x_6_n710), .S(mult_x_6_n711) );
  FA_X1 mult_x_6_U529 ( .A(mult_x_6_n1389), .B(mult_x_6_n711), .CI(
        mult_x_6_n728), .CO(mult_x_6_n708), .S(mult_x_6_n709) );
  FA_X1 mult_x_6_U528 ( .A(mult_x_6_n1421), .B(mult_x_6_n709), .CI(
        mult_x_6_n726), .CO(mult_x_6_n706), .S(mult_x_6_n707) );
  HA_X1 mult_x_6_U527 ( .A(mult_x_6_n724), .B(mult_x_6_n1132), .CO(
        mult_x_6_n704), .S(mult_x_6_n705) );
  FA_X1 mult_x_6_U526 ( .A(mult_x_6_n1164), .B(mult_x_6_n705), .CI(
        mult_x_6_n722), .CO(mult_x_6_n702), .S(mult_x_6_n703) );
  FA_X1 mult_x_6_U525 ( .A(mult_x_6_n1196), .B(mult_x_6_n703), .CI(
        mult_x_6_n720), .CO(mult_x_6_n700), .S(mult_x_6_n701) );
  FA_X1 mult_x_6_U524 ( .A(mult_x_6_n1228), .B(mult_x_6_n701), .CI(
        mult_x_6_n718), .CO(mult_x_6_n698), .S(mult_x_6_n699) );
  FA_X1 mult_x_6_U523 ( .A(mult_x_6_n1260), .B(mult_x_6_n699), .CI(
        mult_x_6_n716), .CO(mult_x_6_n696), .S(mult_x_6_n697) );
  HA_X1 mult_x_6_U517 ( .A(mult_x_6_n704), .B(mult_x_6_n1131), .CO(
        mult_x_6_n684), .S(mult_x_6_n685) );
  FA_X1 mult_x_6_U516 ( .A(mult_x_6_n1163), .B(mult_x_6_n685), .CI(
        mult_x_6_n702), .CO(mult_x_6_n682), .S(mult_x_6_n683) );
  FA_X1 mult_x_6_U515 ( .A(mult_x_6_n1195), .B(mult_x_6_n683), .CI(
        mult_x_6_n700), .CO(mult_x_6_n680), .S(mult_x_6_n681) );
  FA_X1 mult_x_6_U514 ( .A(mult_x_6_n1227), .B(mult_x_6_n681), .CI(
        mult_x_6_n698), .CO(mult_x_6_n678), .S(mult_x_6_n679) );
  FA_X1 mult_x_6_U513 ( .A(mult_x_6_n1259), .B(mult_x_6_n679), .CI(
        mult_x_6_n696), .CO(mult_x_6_n676), .S(mult_x_6_n677) );
  HA_X1 mult_x_6_U507 ( .A(mult_x_6_n684), .B(mult_x_6_n1130), .CO(
        mult_x_6_n664), .S(mult_x_6_n665) );
  FA_X1 mult_x_6_U506 ( .A(mult_x_6_n1162), .B(mult_x_6_n665), .CI(
        mult_x_6_n682), .CO(mult_x_6_n662), .S(mult_x_6_n663) );
  FA_X1 mult_x_6_U505 ( .A(mult_x_6_n1194), .B(mult_x_6_n663), .CI(
        mult_x_6_n680), .CO(mult_x_6_n660), .S(mult_x_6_n661) );
  FA_X1 mult_x_6_U504 ( .A(mult_x_6_n1226), .B(mult_x_6_n661), .CI(
        mult_x_6_n678), .CO(mult_x_6_n658), .S(mult_x_6_n659) );
  FA_X1 mult_x_6_U503 ( .A(mult_x_6_n1258), .B(mult_x_6_n659), .CI(
        mult_x_6_n676), .CO(mult_x_6_n656), .S(mult_x_6_n657) );
  FA_X1 mult_x_6_U502 ( .A(mult_x_6_n1290), .B(mult_x_6_n657), .CI(
        mult_x_6_n674), .CO(mult_x_6_n654), .S(mult_x_6_n655) );
  FA_X1 mult_x_6_U501 ( .A(mult_x_6_n1322), .B(mult_x_6_n655), .CI(
        mult_x_6_n672), .CO(mult_x_6_n652), .S(mult_x_6_n653) );
  FA_X1 mult_x_6_U500 ( .A(mult_x_6_n1354), .B(mult_x_6_n653), .CI(
        mult_x_6_n670), .CO(mult_x_6_n650), .S(mult_x_6_n651) );
  FA_X1 mult_x_6_U498 ( .A(mult_x_6_n1418), .B(mult_x_6_n649), .CI(
        mult_x_6_n666), .CO(mult_x_6_n646), .S(mult_x_6_n647) );
  FA_X1 mult_x_6_U495 ( .A(mult_x_6_n645), .B(mult_x_6_n1129), .CI(
        mult_x_6_n1161), .CO(mult_x_6_n643), .S(mult_x_6_n644) );
  FA_X1 mult_x_6_U494 ( .A(mult_x_6_n644), .B(mult_x_6_n662), .CI(
        mult_x_6_n1193), .CO(mult_x_6_n641), .S(mult_x_6_n642) );
  FA_X1 mult_x_6_U493 ( .A(mult_x_6_n642), .B(mult_x_6_n660), .CI(
        mult_x_6_n1225), .CO(mult_x_6_n639), .S(mult_x_6_n640) );
  FA_X1 mult_x_6_U492 ( .A(mult_x_6_n640), .B(mult_x_6_n658), .CI(
        mult_x_6_n1257), .CO(mult_x_6_n637), .S(mult_x_6_n638) );
  FA_X1 mult_x_6_U491 ( .A(mult_x_6_n638), .B(mult_x_6_n656), .CI(
        mult_x_6_n1289), .CO(mult_x_6_n635), .S(mult_x_6_n636) );
  FA_X1 mult_x_6_U490 ( .A(mult_x_6_n636), .B(mult_x_6_n654), .CI(
        mult_x_6_n1321), .CO(mult_x_6_n633), .S(mult_x_6_n634) );
  FA_X1 mult_x_6_U489 ( .A(mult_x_6_n634), .B(mult_x_6_n652), .CI(
        mult_x_6_n1353), .CO(mult_x_6_n631), .S(mult_x_6_n632) );
  FA_X1 mult_x_6_U488 ( .A(mult_x_6_n632), .B(mult_x_6_n650), .CI(
        mult_x_6_n1385), .CO(mult_x_6_n629), .S(mult_x_6_n630) );
  FA_X1 mult_x_6_U487 ( .A(mult_x_6_n630), .B(mult_x_6_n648), .CI(
        mult_x_6_n1417), .CO(mult_x_6_n627), .S(mult_x_6_n628) );
  FA_X1 mult_x_6_U485 ( .A(mult_x_6_n1128), .B(n2165), .CI(mult_x_6_n1160), 
        .CO(mult_x_6_n624), .S(mult_x_6_n625) );
  FA_X1 mult_x_6_U484 ( .A(mult_x_6_n625), .B(mult_x_6_n643), .CI(
        mult_x_6_n641), .CO(mult_x_6_n622), .S(mult_x_6_n623) );
  FA_X1 mult_x_6_U483 ( .A(mult_x_6_n623), .B(mult_x_6_n1192), .CI(
        mult_x_6_n1224), .CO(mult_x_6_n620), .S(mult_x_6_n621) );
  FA_X1 mult_x_6_U482 ( .A(mult_x_6_n621), .B(mult_x_6_n639), .CI(
        mult_x_6_n637), .CO(mult_x_6_n618), .S(mult_x_6_n619) );
  FA_X1 mult_x_6_U481 ( .A(mult_x_6_n619), .B(mult_x_6_n1256), .CI(
        mult_x_6_n1288), .CO(mult_x_6_n616), .S(mult_x_6_n617) );
  FA_X1 mult_x_6_U480 ( .A(mult_x_6_n617), .B(mult_x_6_n635), .CI(
        mult_x_6_n633), .CO(mult_x_6_n614), .S(mult_x_6_n615) );
  FA_X1 mult_x_6_U479 ( .A(mult_x_6_n615), .B(mult_x_6_n1320), .CI(
        mult_x_6_n1352), .CO(mult_x_6_n612), .S(mult_x_6_n613) );
  FA_X1 mult_x_6_U478 ( .A(mult_x_6_n613), .B(mult_x_6_n631), .CI(
        mult_x_6_n629), .CO(mult_x_6_n610), .S(mult_x_6_n611) );
  FA_X1 mult_x_6_U477 ( .A(mult_x_6_n611), .B(mult_x_6_n1384), .CI(
        mult_x_6_n1416), .CO(mult_x_6_n608), .S(mult_x_6_n609) );
  FA_X1 mult_x_6_U475 ( .A(mult_x_6_n1127), .B(n2165), .CI(mult_x_6_n624), 
        .CO(mult_x_6_n604), .S(mult_x_6_n605) );
  FA_X1 mult_x_6_U474 ( .A(mult_x_6_n605), .B(mult_x_6_n1159), .CI(
        mult_x_6_n622), .CO(mult_x_6_n602), .S(mult_x_6_n603) );
  FA_X1 mult_x_6_U473 ( .A(mult_x_6_n603), .B(mult_x_6_n1191), .CI(
        mult_x_6_n620), .CO(mult_x_6_n600), .S(mult_x_6_n601) );
  FA_X1 mult_x_6_U472 ( .A(mult_x_6_n601), .B(mult_x_6_n1223), .CI(
        mult_x_6_n618), .CO(mult_x_6_n598), .S(mult_x_6_n599) );
  FA_X1 mult_x_6_U471 ( .A(mult_x_6_n599), .B(mult_x_6_n1255), .CI(
        mult_x_6_n1287), .CO(mult_x_6_n596), .S(mult_x_6_n597) );
  FA_X1 mult_x_6_U470 ( .A(mult_x_6_n597), .B(mult_x_6_n616), .CI(
        mult_x_6_n614), .CO(mult_x_6_n594), .S(mult_x_6_n595) );
  FA_X1 mult_x_6_U469 ( .A(mult_x_6_n595), .B(mult_x_6_n1319), .CI(
        mult_x_6_n1351), .CO(mult_x_6_n592), .S(mult_x_6_n593) );
  FA_X1 mult_x_6_U468 ( .A(mult_x_6_n593), .B(mult_x_6_n612), .CI(
        mult_x_6_n610), .CO(mult_x_6_n590), .S(mult_x_6_n591) );
  FA_X1 mult_x_6_U466 ( .A(mult_x_6_n606), .B(mult_x_6_n1414), .CI(
        mult_x_6_n1126), .CO(mult_x_6_n586), .S(mult_x_6_n587) );
  FA_X1 mult_x_6_U465 ( .A(mult_x_6_n604), .B(mult_x_6_n587), .CI(
        mult_x_6_n1158), .CO(mult_x_6_n584), .S(mult_x_6_n585) );
  FA_X1 mult_x_6_U464 ( .A(mult_x_6_n602), .B(mult_x_6_n585), .CI(
        mult_x_6_n1190), .CO(mult_x_6_n582), .S(mult_x_6_n583) );
  FA_X1 mult_x_6_U463 ( .A(mult_x_6_n600), .B(mult_x_6_n583), .CI(
        mult_x_6_n1222), .CO(mult_x_6_n580), .S(mult_x_6_n581) );
  FA_X1 mult_x_6_U462 ( .A(mult_x_6_n1254), .B(mult_x_6_n581), .CI(
        mult_x_6_n598), .CO(mult_x_6_n578), .S(mult_x_6_n579) );
  FA_X1 mult_x_6_U461 ( .A(mult_x_6_n596), .B(mult_x_6_n579), .CI(
        mult_x_6_n1286), .CO(mult_x_6_n576), .S(mult_x_6_n577) );
  FA_X1 mult_x_6_U460 ( .A(mult_x_6_n1318), .B(mult_x_6_n577), .CI(
        mult_x_6_n594), .CO(mult_x_6_n574), .S(mult_x_6_n575) );
  FA_X1 mult_x_6_U459 ( .A(mult_x_6_n592), .B(mult_x_6_n575), .CI(
        mult_x_6_n1350), .CO(mult_x_6_n572), .S(mult_x_6_n573) );
  FA_X1 mult_x_6_U458 ( .A(mult_x_6_n1382), .B(mult_x_6_n573), .CI(
        mult_x_6_n590), .CO(mult_x_6_n570), .S(mult_x_6_n571) );
  FA_X1 mult_x_6_U456 ( .A(n2160), .B(mult_x_6_n586), .CI(mult_x_6_n1157), 
        .CO(mult_x_6_n567), .S(mult_x_6_n568) );
  FA_X1 mult_x_6_U455 ( .A(mult_x_6_n568), .B(mult_x_6_n584), .CI(
        mult_x_6_n1189), .CO(mult_x_6_n565), .S(mult_x_6_n566) );
  FA_X1 mult_x_6_U454 ( .A(mult_x_6_n566), .B(mult_x_6_n582), .CI(
        mult_x_6_n1221), .CO(mult_x_6_n563), .S(mult_x_6_n564) );
  FA_X1 mult_x_6_U453 ( .A(mult_x_6_n564), .B(mult_x_6_n580), .CI(
        mult_x_6_n1253), .CO(mult_x_6_n561), .S(mult_x_6_n562) );
  FA_X1 mult_x_6_U452 ( .A(mult_x_6_n562), .B(mult_x_6_n578), .CI(
        mult_x_6_n1285), .CO(mult_x_6_n559), .S(mult_x_6_n560) );
  FA_X1 mult_x_6_U451 ( .A(mult_x_6_n560), .B(mult_x_6_n576), .CI(
        mult_x_6_n1317), .CO(mult_x_6_n557), .S(mult_x_6_n558) );
  FA_X1 mult_x_6_U450 ( .A(mult_x_6_n558), .B(mult_x_6_n574), .CI(
        mult_x_6_n1349), .CO(mult_x_6_n555), .S(mult_x_6_n556) );
  FA_X1 mult_x_6_U449 ( .A(mult_x_6_n556), .B(mult_x_6_n572), .CI(
        mult_x_6_n1381), .CO(mult_x_6_n553), .S(mult_x_6_n554) );
  FA_X1 mult_x_6_U447 ( .A(mult_x_6_n1125), .B(n2160), .CI(mult_x_6_n1156), 
        .CO(mult_x_6_n549), .S(mult_x_6_n550) );
  FA_X1 mult_x_6_U446 ( .A(mult_x_6_n550), .B(mult_x_6_n567), .CI(
        mult_x_6_n565), .CO(mult_x_6_n547), .S(mult_x_6_n548) );
  FA_X1 mult_x_6_U445 ( .A(mult_x_6_n548), .B(mult_x_6_n1188), .CI(
        mult_x_6_n563), .CO(mult_x_6_n545), .S(mult_x_6_n546) );
  FA_X1 mult_x_6_U444 ( .A(mult_x_6_n546), .B(mult_x_6_n1220), .CI(
        mult_x_6_n1252), .CO(mult_x_6_n543), .S(mult_x_6_n544) );
  FA_X1 mult_x_6_U443 ( .A(mult_x_6_n544), .B(mult_x_6_n561), .CI(
        mult_x_6_n559), .CO(mult_x_6_n541), .S(mult_x_6_n542) );
  FA_X1 mult_x_6_U442 ( .A(mult_x_6_n542), .B(mult_x_6_n1284), .CI(
        mult_x_6_n1316), .CO(mult_x_6_n539), .S(mult_x_6_n540) );
  FA_X1 mult_x_6_U441 ( .A(mult_x_6_n540), .B(mult_x_6_n557), .CI(
        mult_x_6_n555), .CO(mult_x_6_n537), .S(mult_x_6_n538) );
  FA_X1 mult_x_6_U440 ( .A(mult_x_6_n1380), .B(mult_x_6_n1348), .CI(
        mult_x_6_n538), .CO(mult_x_6_n535), .S(mult_x_6_n536) );
  FA_X1 mult_x_6_U439 ( .A(mult_x_6_n551), .B(mult_x_6_n1379), .CI(
        mult_x_6_n1124), .CO(mult_x_6_n503), .S(mult_x_6_n534) );
  FA_X1 mult_x_6_U438 ( .A(mult_x_6_n549), .B(mult_x_6_n534), .CI(
        mult_x_6_n1155), .CO(mult_x_6_n532), .S(mult_x_6_n533) );
  FA_X1 mult_x_6_U437 ( .A(mult_x_6_n547), .B(mult_x_6_n533), .CI(
        mult_x_6_n1187), .CO(mult_x_6_n530), .S(mult_x_6_n531) );
  FA_X1 mult_x_6_U436 ( .A(mult_x_6_n1219), .B(mult_x_6_n531), .CI(
        mult_x_6_n545), .CO(mult_x_6_n528), .S(mult_x_6_n529) );
  FA_X1 mult_x_6_U435 ( .A(mult_x_6_n543), .B(mult_x_6_n529), .CI(
        mult_x_6_n1251), .CO(mult_x_6_n526), .S(mult_x_6_n527) );
  FA_X1 mult_x_6_U434 ( .A(mult_x_6_n1283), .B(mult_x_6_n527), .CI(
        mult_x_6_n541), .CO(mult_x_6_n524), .S(mult_x_6_n525) );
  FA_X1 mult_x_6_U433 ( .A(mult_x_6_n539), .B(mult_x_6_n525), .CI(
        mult_x_6_n1315), .CO(mult_x_6_n522), .S(mult_x_6_n523) );
  FA_X1 mult_x_6_U432 ( .A(mult_x_6_n1347), .B(mult_x_6_n523), .CI(
        mult_x_6_n537), .CO(mult_x_6_n520), .S(mult_x_6_n521) );
  FA_X1 mult_x_6_U430 ( .A(n2166), .B(mult_x_6_n1123), .CI(mult_x_6_n1154), 
        .CO(mult_x_6_n517), .S(mult_x_6_n518) );
  FA_X1 mult_x_6_U429 ( .A(mult_x_6_n518), .B(mult_x_6_n532), .CI(
        mult_x_6_n1186), .CO(mult_x_6_n515), .S(mult_x_6_n516) );
  FA_X1 mult_x_6_U428 ( .A(mult_x_6_n516), .B(mult_x_6_n530), .CI(
        mult_x_6_n1218), .CO(mult_x_6_n513), .S(mult_x_6_n514) );
  FA_X1 mult_x_6_U427 ( .A(mult_x_6_n514), .B(mult_x_6_n528), .CI(
        mult_x_6_n1250), .CO(mult_x_6_n511), .S(mult_x_6_n512) );
  FA_X1 mult_x_6_U426 ( .A(mult_x_6_n512), .B(mult_x_6_n526), .CI(
        mult_x_6_n1282), .CO(mult_x_6_n509), .S(mult_x_6_n510) );
  FA_X1 mult_x_6_U425 ( .A(mult_x_6_n510), .B(mult_x_6_n524), .CI(
        mult_x_6_n1314), .CO(mult_x_6_n507), .S(mult_x_6_n508) );
  FA_X1 mult_x_6_U424 ( .A(mult_x_6_n508), .B(mult_x_6_n522), .CI(
        mult_x_6_n1346), .CO(mult_x_6_n505), .S(mult_x_6_n506) );
  FA_X1 mult_x_6_U422 ( .A(mult_x_6_n1122), .B(n2166), .CI(mult_x_6_n517), 
        .CO(mult_x_6_n501), .S(mult_x_6_n502) );
  FA_X1 mult_x_6_U421 ( .A(mult_x_6_n502), .B(mult_x_6_n1153), .CI(
        mult_x_6_n515), .CO(mult_x_6_n499), .S(mult_x_6_n500) );
  FA_X1 mult_x_6_U420 ( .A(mult_x_6_n500), .B(mult_x_6_n1185), .CI(
        mult_x_6_n1217), .CO(mult_x_6_n497), .S(mult_x_6_n498) );
  FA_X1 mult_x_6_U419 ( .A(mult_x_6_n498), .B(mult_x_6_n513), .CI(
        mult_x_6_n511), .CO(mult_x_6_n495), .S(mult_x_6_n496) );
  FA_X1 mult_x_6_U418 ( .A(mult_x_6_n496), .B(mult_x_6_n1249), .CI(
        mult_x_6_n1281), .CO(mult_x_6_n493), .S(mult_x_6_n494) );
  FA_X1 mult_x_6_U417 ( .A(mult_x_6_n494), .B(mult_x_6_n509), .CI(
        mult_x_6_n507), .CO(mult_x_6_n491), .S(mult_x_6_n492) );
  FA_X1 mult_x_6_U416 ( .A(mult_x_6_n1345), .B(mult_x_6_n1313), .CI(
        mult_x_6_n492), .CO(mult_x_6_n489), .S(mult_x_6_n490) );
  FA_X1 mult_x_6_U415 ( .A(mult_x_6_n503), .B(mult_x_6_n1344), .CI(
        mult_x_6_n1121), .CO(mult_x_6_n487), .S(mult_x_6_n488) );
  FA_X1 mult_x_6_U414 ( .A(mult_x_6_n501), .B(mult_x_6_n488), .CI(
        mult_x_6_n1152), .CO(mult_x_6_n485), .S(mult_x_6_n486) );
  FA_X1 mult_x_6_U413 ( .A(mult_x_6_n1184), .B(mult_x_6_n486), .CI(
        mult_x_6_n499), .CO(mult_x_6_n483), .S(mult_x_6_n484) );
  FA_X1 mult_x_6_U412 ( .A(mult_x_6_n497), .B(mult_x_6_n484), .CI(
        mult_x_6_n1216), .CO(mult_x_6_n481), .S(mult_x_6_n482) );
  FA_X1 mult_x_6_U411 ( .A(mult_x_6_n1248), .B(mult_x_6_n482), .CI(
        mult_x_6_n495), .CO(mult_x_6_n479), .S(mult_x_6_n480) );
  FA_X1 mult_x_6_U410 ( .A(mult_x_6_n493), .B(mult_x_6_n480), .CI(
        mult_x_6_n1280), .CO(mult_x_6_n477), .S(mult_x_6_n478) );
  FA_X1 mult_x_6_U409 ( .A(mult_x_6_n1312), .B(mult_x_6_n478), .CI(
        mult_x_6_n491), .CO(mult_x_6_n475), .S(mult_x_6_n476) );
  FA_X1 mult_x_6_U407 ( .A(n2161), .B(mult_x_6_n487), .CI(mult_x_6_n1151), 
        .CO(mult_x_6_n472), .S(mult_x_6_n473) );
  FA_X1 mult_x_6_U406 ( .A(mult_x_6_n473), .B(mult_x_6_n485), .CI(
        mult_x_6_n1183), .CO(mult_x_6_n470), .S(mult_x_6_n471) );
  FA_X1 mult_x_6_U405 ( .A(mult_x_6_n471), .B(mult_x_6_n483), .CI(
        mult_x_6_n1215), .CO(mult_x_6_n468), .S(mult_x_6_n469) );
  FA_X1 mult_x_6_U404 ( .A(mult_x_6_n469), .B(mult_x_6_n481), .CI(
        mult_x_6_n1247), .CO(mult_x_6_n466), .S(mult_x_6_n467) );
  FA_X1 mult_x_6_U403 ( .A(mult_x_6_n467), .B(mult_x_6_n479), .CI(
        mult_x_6_n1279), .CO(mult_x_6_n464), .S(mult_x_6_n465) );
  FA_X1 mult_x_6_U402 ( .A(mult_x_6_n465), .B(mult_x_6_n477), .CI(
        mult_x_6_n1311), .CO(mult_x_6_n462), .S(mult_x_6_n463) );
  FA_X1 mult_x_6_U400 ( .A(mult_x_6_n1120), .B(n2161), .CI(mult_x_6_n472), 
        .CO(mult_x_6_n458), .S(mult_x_6_n459) );
  FA_X1 mult_x_6_U399 ( .A(mult_x_6_n459), .B(mult_x_6_n1150), .CI(
        mult_x_6_n1182), .CO(mult_x_6_n456), .S(mult_x_6_n457) );
  FA_X1 mult_x_6_U398 ( .A(mult_x_6_n457), .B(mult_x_6_n470), .CI(
        mult_x_6_n468), .CO(mult_x_6_n454), .S(mult_x_6_n455) );
  FA_X1 mult_x_6_U397 ( .A(mult_x_6_n455), .B(mult_x_6_n1214), .CI(
        mult_x_6_n1246), .CO(mult_x_6_n452), .S(mult_x_6_n453) );
  FA_X1 mult_x_6_U396 ( .A(mult_x_6_n453), .B(mult_x_6_n466), .CI(
        mult_x_6_n464), .CO(mult_x_6_n450), .S(mult_x_6_n451) );
  FA_X1 mult_x_6_U395 ( .A(mult_x_6_n1310), .B(mult_x_6_n1278), .CI(
        mult_x_6_n451), .CO(mult_x_6_n448), .S(mult_x_6_n449) );
  FA_X1 mult_x_6_U394 ( .A(mult_x_6_n460), .B(mult_x_6_n1309), .CI(
        mult_x_6_n1119), .CO(mult_x_6_n424), .S(mult_x_6_n447) );
  FA_X1 mult_x_6_U393 ( .A(mult_x_6_n1149), .B(mult_x_6_n447), .CI(
        mult_x_6_n458), .CO(mult_x_6_n445), .S(mult_x_6_n446) );
  FA_X1 mult_x_6_U392 ( .A(mult_x_6_n456), .B(mult_x_6_n446), .CI(
        mult_x_6_n1181), .CO(mult_x_6_n443), .S(mult_x_6_n444) );
  FA_X1 mult_x_6_U391 ( .A(mult_x_6_n1213), .B(mult_x_6_n444), .CI(
        mult_x_6_n454), .CO(mult_x_6_n441), .S(mult_x_6_n442) );
  FA_X1 mult_x_6_U390 ( .A(mult_x_6_n452), .B(mult_x_6_n442), .CI(
        mult_x_6_n1245), .CO(mult_x_6_n439), .S(mult_x_6_n440) );
  FA_X1 mult_x_6_U389 ( .A(mult_x_6_n1277), .B(mult_x_6_n440), .CI(
        mult_x_6_n450), .CO(mult_x_6_n437), .S(mult_x_6_n438) );
  FA_X1 mult_x_6_U387 ( .A(n2167), .B(mult_x_6_n1118), .CI(mult_x_6_n1148), 
        .CO(mult_x_6_n434), .S(mult_x_6_n435) );
  FA_X1 mult_x_6_U386 ( .A(mult_x_6_n435), .B(mult_x_6_n445), .CI(
        mult_x_6_n1180), .CO(mult_x_6_n432), .S(mult_x_6_n433) );
  FA_X1 mult_x_6_U385 ( .A(mult_x_6_n433), .B(mult_x_6_n443), .CI(
        mult_x_6_n1212), .CO(mult_x_6_n430), .S(mult_x_6_n431) );
  FA_X1 mult_x_6_U384 ( .A(mult_x_6_n431), .B(mult_x_6_n441), .CI(
        mult_x_6_n1244), .CO(mult_x_6_n428), .S(mult_x_6_n429) );
  FA_X1 mult_x_6_U383 ( .A(mult_x_6_n429), .B(mult_x_6_n439), .CI(
        mult_x_6_n1276), .CO(mult_x_6_n426), .S(mult_x_6_n427) );
  FA_X1 mult_x_6_U381 ( .A(mult_x_6_n1117), .B(n2167), .CI(mult_x_6_n1147), 
        .CO(mult_x_6_n422), .S(mult_x_6_n423) );
  FA_X1 mult_x_6_U380 ( .A(mult_x_6_n423), .B(mult_x_6_n434), .CI(
        mult_x_6_n432), .CO(mult_x_6_n420), .S(mult_x_6_n421) );
  FA_X1 mult_x_6_U379 ( .A(mult_x_6_n421), .B(mult_x_6_n1179), .CI(
        mult_x_6_n1211), .CO(mult_x_6_n418), .S(mult_x_6_n419) );
  FA_X1 mult_x_6_U378 ( .A(mult_x_6_n419), .B(mult_x_6_n430), .CI(
        mult_x_6_n428), .CO(mult_x_6_n416), .S(mult_x_6_n417) );
  FA_X1 mult_x_6_U377 ( .A(mult_x_6_n1275), .B(mult_x_6_n1243), .CI(
        mult_x_6_n417), .CO(mult_x_6_n414), .S(mult_x_6_n415) );
  FA_X1 mult_x_6_U376 ( .A(mult_x_6_n424), .B(mult_x_6_n1274), .CI(
        mult_x_6_n1116), .CO(mult_x_6_n412), .S(mult_x_6_n413) );
  FA_X1 mult_x_6_U375 ( .A(mult_x_6_n422), .B(mult_x_6_n413), .CI(
        mult_x_6_n1146), .CO(mult_x_6_n410), .S(mult_x_6_n411) );
  FA_X1 mult_x_6_U374 ( .A(mult_x_6_n1178), .B(mult_x_6_n411), .CI(
        mult_x_6_n420), .CO(mult_x_6_n408), .S(mult_x_6_n409) );
  FA_X1 mult_x_6_U373 ( .A(mult_x_6_n418), .B(mult_x_6_n409), .CI(
        mult_x_6_n1210), .CO(mult_x_6_n406), .S(mult_x_6_n407) );
  FA_X1 mult_x_6_U372 ( .A(mult_x_6_n1242), .B(mult_x_6_n407), .CI(
        mult_x_6_n416), .CO(mult_x_6_n404), .S(mult_x_6_n405) );
  FA_X1 mult_x_6_U370 ( .A(n2162), .B(mult_x_6_n412), .CI(mult_x_6_n1145), 
        .CO(mult_x_6_n401), .S(mult_x_6_n402) );
  FA_X1 mult_x_6_U369 ( .A(mult_x_6_n402), .B(mult_x_6_n410), .CI(
        mult_x_6_n1177), .CO(mult_x_6_n399), .S(mult_x_6_n400) );
  FA_X1 mult_x_6_U368 ( .A(mult_x_6_n400), .B(mult_x_6_n408), .CI(
        mult_x_6_n1209), .CO(mult_x_6_n397), .S(mult_x_6_n398) );
  FA_X1 mult_x_6_U367 ( .A(mult_x_6_n398), .B(mult_x_6_n406), .CI(
        mult_x_6_n1241), .CO(mult_x_6_n395), .S(mult_x_6_n396) );
  FA_X1 mult_x_6_U365 ( .A(mult_x_6_n1115), .B(n2162), .CI(mult_x_6_n401), 
        .CO(mult_x_6_n391), .S(mult_x_6_n392) );
  FA_X1 mult_x_6_U364 ( .A(mult_x_6_n392), .B(mult_x_6_n1144), .CI(
        mult_x_6_n1176), .CO(mult_x_6_n389), .S(mult_x_6_n390) );
  FA_X1 mult_x_6_U363 ( .A(mult_x_6_n390), .B(mult_x_6_n399), .CI(
        mult_x_6_n397), .CO(mult_x_6_n387), .S(mult_x_6_n388) );
  FA_X1 mult_x_6_U362 ( .A(mult_x_6_n1240), .B(mult_x_6_n1208), .CI(
        mult_x_6_n388), .CO(mult_x_6_n385), .S(mult_x_6_n386) );
  FA_X1 mult_x_6_U361 ( .A(mult_x_6_n393), .B(mult_x_6_n1239), .CI(
        mult_x_6_n1114), .CO(mult_x_6_n369), .S(mult_x_6_n384) );
  FA_X1 mult_x_6_U360 ( .A(mult_x_6_n1143), .B(mult_x_6_n384), .CI(
        mult_x_6_n391), .CO(mult_x_6_n382), .S(mult_x_6_n383) );
  FA_X1 mult_x_6_U359 ( .A(mult_x_6_n389), .B(mult_x_6_n383), .CI(
        mult_x_6_n1175), .CO(mult_x_6_n380), .S(mult_x_6_n381) );
  FA_X1 mult_x_6_U358 ( .A(mult_x_6_n1207), .B(mult_x_6_n381), .CI(
        mult_x_6_n387), .CO(mult_x_6_n378), .S(mult_x_6_n379) );
  FA_X1 mult_x_6_U356 ( .A(n2168), .B(mult_x_6_n1113), .CI(mult_x_6_n1142), 
        .CO(mult_x_6_n375), .S(mult_x_6_n376) );
  FA_X1 mult_x_6_U355 ( .A(mult_x_6_n376), .B(mult_x_6_n382), .CI(
        mult_x_6_n1174), .CO(mult_x_6_n373), .S(mult_x_6_n374) );
  FA_X1 mult_x_6_U354 ( .A(mult_x_6_n374), .B(mult_x_6_n380), .CI(
        mult_x_6_n1206), .CO(mult_x_6_n371), .S(mult_x_6_n372) );
  FA_X1 mult_x_6_U352 ( .A(mult_x_6_n1112), .B(n2168), .CI(mult_x_6_n1141), 
        .CO(mult_x_6_n367), .S(mult_x_6_n368) );
  FA_X1 mult_x_6_U351 ( .A(mult_x_6_n368), .B(mult_x_6_n375), .CI(
        mult_x_6_n373), .CO(mult_x_6_n365), .S(mult_x_6_n366) );
  FA_X1 mult_x_6_U350 ( .A(mult_x_6_n1205), .B(mult_x_6_n1173), .CI(
        mult_x_6_n366), .CO(mult_x_6_n363), .S(mult_x_6_n364) );
  FA_X1 mult_x_6_U349 ( .A(mult_x_6_n369), .B(mult_x_6_n1204), .CI(
        mult_x_6_n1111), .CO(mult_x_6_n361), .S(mult_x_6_n362) );
  FA_X1 mult_x_6_U348 ( .A(mult_x_6_n367), .B(mult_x_6_n362), .CI(
        mult_x_6_n1140), .CO(mult_x_6_n359), .S(mult_x_6_n360) );
  FA_X1 mult_x_6_U347 ( .A(mult_x_6_n1172), .B(mult_x_6_n360), .CI(
        mult_x_6_n365), .CO(mult_x_6_n357), .S(mult_x_6_n358) );
  FA_X1 mult_x_6_U345 ( .A(n2163), .B(mult_x_6_n361), .CI(mult_x_6_n1139), 
        .CO(mult_x_6_n354), .S(mult_x_6_n355) );
  FA_X1 mult_x_6_U344 ( .A(mult_x_6_n355), .B(mult_x_6_n359), .CI(
        mult_x_6_n1171), .CO(mult_x_6_n352), .S(mult_x_6_n353) );
  FA_X1 mult_x_6_U342 ( .A(mult_x_6_n1110), .B(n2163), .CI(mult_x_6_n354), 
        .CO(mult_x_6_n348), .S(mult_x_6_n349) );
  FA_X1 mult_x_6_U341 ( .A(mult_x_6_n1170), .B(mult_x_6_n1138), .CI(
        mult_x_6_n349), .CO(mult_x_6_n346), .S(mult_x_6_n347) );
  FA_X1 mult_x_6_U340 ( .A(mult_x_6_n350), .B(mult_x_6_n1169), .CI(
        mult_x_6_n1109), .CO(mult_x_6_n338), .S(mult_x_6_n345) );
  FA_X1 mult_x_6_U339 ( .A(mult_x_6_n1137), .B(mult_x_6_n345), .CI(
        mult_x_6_n348), .CO(mult_x_6_n343), .S(mult_x_6_n344) );
  FA_X1 mult_x_6_U337 ( .A(n2169), .B(mult_x_6_n1108), .CI(mult_x_6_n1136), 
        .CO(mult_x_6_n340), .S(mult_x_6_n341) );
  FA_X1 mult_x_6_U335 ( .A(mult_x_6_n1107), .B(n2169), .CI(mult_x_6_n1135), 
        .CO(mult_x_6_n336), .S(mult_x_6_n337) );
  FA_X1 mult_x_6_U334 ( .A(mult_x_6_n338), .B(mult_x_6_n1134), .CI(
        mult_x_6_n1106), .CO(mult_x_6_n334), .S(mult_x_6_n335) );
  HA_X1 mult_x_6_U331 ( .A(mult_x_6_n1483), .B(mul_operand_a_q[2]), .CO(
        mult_x_6_n330), .S(mult_result_w[0]) );
  FA_X1 mult_x_6_U327 ( .A(mult_x_6_n1479), .B(mult_x_6_n993), .CI(
        mult_x_6_n327), .CO(mult_x_6_n326), .S(mult_result_w[4]) );
  FA_X1 mult_x_6_U326 ( .A(mult_x_6_n1478), .B(mult_x_6_n991), .CI(
        mult_x_6_n326), .CO(mult_x_6_n325), .S(mult_result_w[5]) );
  FA_X1 mult_x_6_U324 ( .A(mult_x_6_n1476), .B(mult_x_6_n983), .CI(
        mult_x_6_n324), .CO(mult_x_6_n323), .S(mult_result_w[7]) );
  FA_X1 mult_x_6_U314 ( .A(mult_x_6_n1466), .B(mult_x_6_n907), .CI(
        mult_x_6_n314), .CO(mult_x_6_n313), .S(mult_result_w[17]) );
  FA_X1 mult_x_6_U313 ( .A(mult_x_6_n1465), .B(mult_x_6_n895), .CI(
        mult_x_6_n313), .CO(mult_x_6_n312), .S(mult_result_w[18]) );
  FA_X1 mult_x_6_U308 ( .A(mult_x_6_n1460), .B(mult_x_6_n829), .CI(
        mult_x_6_n308), .CO(mult_x_6_n307), .S(mult_result_w[23]) );
  FA_X1 mult_x_6_U300 ( .A(mult_x_6_n1452), .B(mult_x_6_n687), .CI(
        mult_x_6_n300), .CO(mult_x_6_n299), .S(mult_result_w[31]) );
  OR2_X1 DP_OP_56J3_124_887_U34 ( .A1(n1028), .A2(C1_Z_0), .ZN(
        DP_OP_56J3_124_887_n32) );
  XNOR2_X1 DP_OP_56J3_124_887_U33 ( .A(n1028), .B(C1_Z_0), .ZN(C21_DATA3_0) );
  FA_X1 DP_OP_56J3_124_887_U32 ( .A(n1029), .B(C1_Z_1), .CI(
        DP_OP_56J3_124_887_n32), .CO(DP_OP_56J3_124_887_n31), .S(C21_DATA3_1)
         );
  FA_X1 DP_OP_56J3_124_887_U31 ( .A(n1040), .B(C1_Z_2), .CI(
        DP_OP_56J3_124_887_n31), .CO(DP_OP_56J3_124_887_n30), .S(C21_DATA3_2)
         );
  FA_X1 DP_OP_56J3_124_887_U30 ( .A(n1051), .B(C1_Z_3), .CI(
        DP_OP_56J3_124_887_n30), .CO(DP_OP_56J3_124_887_n29), .S(C21_DATA3_3)
         );
  FA_X1 DP_OP_56J3_124_887_U29 ( .A(n1053), .B(C1_Z_4), .CI(
        DP_OP_56J3_124_887_n29), .CO(DP_OP_56J3_124_887_n28), .S(C21_DATA3_4)
         );
  FA_X1 DP_OP_56J3_124_887_U28 ( .A(n1054), .B(C1_Z_5), .CI(
        DP_OP_56J3_124_887_n28), .CO(DP_OP_56J3_124_887_n27), .S(C21_DATA3_5)
         );
  FA_X1 DP_OP_56J3_124_887_U27 ( .A(n1055), .B(C1_Z_6), .CI(
        DP_OP_56J3_124_887_n27), .CO(DP_OP_56J3_124_887_n26), .S(C21_DATA3_6)
         );
  FA_X1 DP_OP_56J3_124_887_U26 ( .A(n1056), .B(C1_Z_7), .CI(
        DP_OP_56J3_124_887_n26), .CO(DP_OP_56J3_124_887_n25), .S(C21_DATA3_7)
         );
  FA_X1 DP_OP_56J3_124_887_U25 ( .A(n1057), .B(C1_Z_8), .CI(
        DP_OP_56J3_124_887_n25), .CO(DP_OP_56J3_124_887_n24), .S(C21_DATA3_8)
         );
  FA_X1 DP_OP_56J3_124_887_U24 ( .A(n1058), .B(C1_Z_9), .CI(
        DP_OP_56J3_124_887_n24), .CO(DP_OP_56J3_124_887_n23), .S(C21_DATA3_9)
         );
  FA_X1 DP_OP_56J3_124_887_U23 ( .A(n1030), .B(C1_Z_10), .CI(
        DP_OP_56J3_124_887_n23), .CO(DP_OP_56J3_124_887_n22), .S(C21_DATA3_10)
         );
  FA_X1 DP_OP_56J3_124_887_U22 ( .A(n1031), .B(C1_Z_11), .CI(
        DP_OP_56J3_124_887_n22), .CO(DP_OP_56J3_124_887_n21), .S(C21_DATA3_11)
         );
  FA_X1 DP_OP_56J3_124_887_U21 ( .A(n1032), .B(C1_Z_12), .CI(
        DP_OP_56J3_124_887_n21), .CO(DP_OP_56J3_124_887_n20), .S(C21_DATA3_12)
         );
  FA_X1 DP_OP_56J3_124_887_U20 ( .A(n1033), .B(C1_Z_13), .CI(
        DP_OP_56J3_124_887_n20), .CO(DP_OP_56J3_124_887_n19), .S(C21_DATA3_13)
         );
  FA_X1 DP_OP_56J3_124_887_U19 ( .A(n1034), .B(C1_Z_14), .CI(
        DP_OP_56J3_124_887_n19), .CO(DP_OP_56J3_124_887_n18), .S(C21_DATA3_14)
         );
  FA_X1 DP_OP_56J3_124_887_U18 ( .A(n1035), .B(C1_Z_15), .CI(
        DP_OP_56J3_124_887_n18), .CO(DP_OP_56J3_124_887_n17), .S(C21_DATA3_15)
         );
  FA_X1 DP_OP_56J3_124_887_U17 ( .A(n1036), .B(C1_Z_16), .CI(
        DP_OP_56J3_124_887_n17), .CO(DP_OP_56J3_124_887_n16), .S(C21_DATA3_16)
         );
  FA_X1 DP_OP_56J3_124_887_U16 ( .A(n1037), .B(C1_Z_17), .CI(
        DP_OP_56J3_124_887_n16), .CO(DP_OP_56J3_124_887_n15), .S(C21_DATA3_17)
         );
  FA_X1 DP_OP_56J3_124_887_U15 ( .A(n1038), .B(C1_Z_18), .CI(
        DP_OP_56J3_124_887_n15), .CO(DP_OP_56J3_124_887_n14), .S(C21_DATA3_18)
         );
  FA_X1 DP_OP_56J3_124_887_U14 ( .A(n1039), .B(C1_Z_19), .CI(
        DP_OP_56J3_124_887_n14), .CO(DP_OP_56J3_124_887_n13), .S(C21_DATA3_19)
         );
  FA_X1 DP_OP_56J3_124_887_U13 ( .A(n1041), .B(C1_Z_20), .CI(
        DP_OP_56J3_124_887_n13), .CO(DP_OP_56J3_124_887_n12), .S(C21_DATA3_20)
         );
  FA_X1 DP_OP_56J3_124_887_U12 ( .A(n1042), .B(C1_Z_21), .CI(
        DP_OP_56J3_124_887_n12), .CO(DP_OP_56J3_124_887_n11), .S(C21_DATA3_21)
         );
  FA_X1 DP_OP_56J3_124_887_U11 ( .A(n1043), .B(C1_Z_22), .CI(
        DP_OP_56J3_124_887_n11), .CO(DP_OP_56J3_124_887_n10), .S(C21_DATA3_22)
         );
  FA_X1 DP_OP_56J3_124_887_U10 ( .A(n1044), .B(C1_Z_23), .CI(
        DP_OP_56J3_124_887_n10), .CO(DP_OP_56J3_124_887_n9), .S(C21_DATA3_23)
         );
  FA_X1 DP_OP_56J3_124_887_U9 ( .A(n1045), .B(C1_Z_24), .CI(
        DP_OP_56J3_124_887_n9), .CO(DP_OP_56J3_124_887_n8), .S(C21_DATA3_24)
         );
  FA_X1 DP_OP_56J3_124_887_U8 ( .A(n1046), .B(C1_Z_25), .CI(
        DP_OP_56J3_124_887_n8), .CO(DP_OP_56J3_124_887_n7), .S(C21_DATA3_25)
         );
  FA_X1 DP_OP_56J3_124_887_U7 ( .A(n1047), .B(C1_Z_26), .CI(
        DP_OP_56J3_124_887_n7), .CO(DP_OP_56J3_124_887_n6), .S(C21_DATA3_26)
         );
  FA_X1 DP_OP_56J3_124_887_U6 ( .A(n1048), .B(C1_Z_27), .CI(
        DP_OP_56J3_124_887_n6), .CO(DP_OP_56J3_124_887_n5), .S(C21_DATA3_27)
         );
  FA_X1 DP_OP_56J3_124_887_U5 ( .A(n1049), .B(C1_Z_28), .CI(
        DP_OP_56J3_124_887_n5), .CO(DP_OP_56J3_124_887_n4), .S(C21_DATA3_28)
         );
  FA_X1 DP_OP_56J3_124_887_U4 ( .A(n1050), .B(C1_Z_29), .CI(
        DP_OP_56J3_124_887_n4), .CO(DP_OP_56J3_124_887_n3), .S(C21_DATA3_29)
         );
  FA_X1 DP_OP_56J3_124_887_U3 ( .A(n1052), .B(C1_Z_30), .CI(
        DP_OP_56J3_124_887_n3), .CO(DP_OP_56J3_124_887_n2), .S(C21_DATA3_30)
         );
  XOR2_X1 DP_OP_56J3_124_887_U2 ( .A(DP_OP_56J3_124_887_n132), .B(C1_Z_31), 
        .Z(DP_OP_56J3_124_887_n1) );
  SDFF_X1 mul_operand_a_q_reg_2_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[2]), 
        .CK(clk_i), .Q(mul_operand_a_q[2]), .QN(n1025) );
  DFF_X1 mul_operand_b_q_reg_1_ ( .D(N57), .CK(clk_i), .Q(mul_operand_b_q[1]), 
        .QN(n1021) );
  DFF_X1 result_q_reg_30_ ( .D(n447), .CK(clk_i), .Q(result_o[30]) );
  SDFF_X1 mul_operand_b_q_reg_31_ ( .D(1'b0), .SI(n611), .SE(operand_rb_i[31]), 
        .CK(clk_i), .Q(mul_operand_b_q[31]), .QN(n2178) );
  SDFF_X1 mul_operand_a_q_reg_31_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[31]), 
        .CK(clk_i), .Q(mul_operand_a_q[31]) );
  SDFF_X1 mul_operand_a_q_reg_30_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[30]), 
        .CK(clk_i), .Q(mul_operand_a_q[30]) );
  SDFF_X1 mul_operand_a_q_reg_28_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[28]), 
        .CK(clk_i), .Q(mul_operand_a_q[28]) );
  SDFF_X1 mul_operand_a_q_reg_27_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[27]), 
        .CK(clk_i), .Q(mul_operand_a_q[27]) );
  SDFF_X1 mul_operand_a_q_reg_25_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[25]), 
        .CK(clk_i), .Q(mul_operand_a_q[25]) );
  SDFF_X1 mul_operand_a_q_reg_24_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[24]), 
        .CK(clk_i), .Q(mul_operand_a_q[24]) );
  SDFF_X1 mul_operand_a_q_reg_22_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[22]), 
        .CK(clk_i), .Q(mul_operand_a_q[22]) );
  SDFF_X1 mul_operand_a_q_reg_21_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[21]), 
        .CK(clk_i), .Q(mul_operand_a_q[21]) );
  SDFF_X1 mul_operand_a_q_reg_20_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[20]), 
        .CK(clk_i), .Q(mul_operand_a_q[20]) );
  SDFF_X1 mul_operand_a_q_reg_19_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[19]), 
        .CK(clk_i), .Q(mul_operand_a_q[19]) );
  SDFF_X1 mul_operand_a_q_reg_18_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[18]), 
        .CK(clk_i), .Q(mul_operand_a_q[18]) );
  SDFF_X1 mul_operand_a_q_reg_17_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[17]), 
        .CK(clk_i), .Q(mul_operand_a_q[17]) );
  SDFF_X1 mul_operand_a_q_reg_16_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[16]), 
        .CK(clk_i), .Q(mul_operand_a_q[16]) );
  SDFF_X1 mul_operand_a_q_reg_15_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[15]), 
        .CK(clk_i), .Q(mul_operand_a_q[15]) );
  SDFF_X1 mul_operand_a_q_reg_14_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[14]), 
        .CK(clk_i), .Q(mul_operand_a_q[14]) );
  SDFF_X1 mul_operand_a_q_reg_13_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[13]), 
        .CK(clk_i), .Q(mul_operand_a_q[13]) );
  SDFF_X1 mul_operand_a_q_reg_12_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[12]), 
        .CK(clk_i), .Q(mul_operand_a_q[12]) );
  SDFF_X1 mul_operand_a_q_reg_11_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[11]), 
        .CK(clk_i), .Q(mul_operand_a_q[11]) );
  SDFF_X1 mul_operand_a_q_reg_10_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[10]), 
        .CK(clk_i), .Q(mul_operand_a_q[10]) );
  SDFF_X1 mul_operand_a_q_reg_9_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[9]), 
        .CK(clk_i), .Q(mul_operand_a_q[9]) );
  SDFF_X1 mul_operand_a_q_reg_8_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[8]), 
        .CK(clk_i), .Q(mul_operand_a_q[8]), .QN(n348) );
  DFF_X1 ready_q_reg ( .D(N575), .CK(clk_i), .Q(ready_o) );
  DFF_X1 mul_operand_b_q_reg_32_ ( .D(N88), .CK(clk_i), .Q(mul_operand_b_q[32]) );
  DFF_X1 mul_operand_b_q_reg_30_ ( .D(N86), .CK(clk_i), .Q(mul_operand_b_q[30]) );
  DFF_X1 mul_operand_b_q_reg_28_ ( .D(N84), .CK(clk_i), .Q(mul_operand_b_q[28]), .QN(n353) );
  DFF_X1 mul_operand_b_q_reg_26_ ( .D(N82), .CK(clk_i), .Q(mul_operand_b_q[26]), .QN(n354) );
  DFF_X1 mul_operand_b_q_reg_24_ ( .D(N80), .CK(clk_i), .Q(mul_operand_b_q[24]) );
  DFF_X1 mul_operand_b_q_reg_16_ ( .D(N72), .CK(clk_i), .Q(mul_operand_b_q[16]) );
  DFF_X1 mul_operand_b_q_reg_9_ ( .D(N65), .CK(clk_i), .Q(mul_operand_b_q[9])
         );
  DFF_X1 mul_operand_b_q_reg_6_ ( .D(N62), .CK(clk_i), .Q(mul_operand_b_q[6])
         );
  DFF_X1 mul_operand_b_q_reg_5_ ( .D(N61), .CK(clk_i), .Q(mul_operand_b_q[5])
         );
  DFF_X1 mul_operand_b_q_reg_3_ ( .D(N59), .CK(clk_i), .Q(mul_operand_b_q[3])
         );
  DFF_X1 mul_operand_a_q_reg_7_ ( .D(n2534), .CK(clk_i), .Q(mul_operand_a_q[7]) );
  DFF_X1 mul_operand_a_q_reg_4_ ( .D(n2532), .CK(clk_i), .Q(mul_operand_a_q[4]) );
  DFF_X1 mul_operand_a_q_reg_3_ ( .D(n2531), .CK(clk_i), .Q(mul_operand_a_q[3]) );
  DFF_X1 mul_operand_a_q_reg_0_ ( .D(n2529), .CK(clk_i), .Q(mul_operand_a_q[0]), .QN(n2405) );
  DFF_X1 mul_operand_a_q_reg_6_ ( .D(n2533), .CK(clk_i), .Q(mul_operand_a_q[6]) );
  DFF_X1 divisor_q_reg_33_ ( .D(n542), .CK(clk_i), .Q(divisor_q[33]) );
  DFF_X1 divisor_q_reg_45_ ( .D(n530), .CK(clk_i), .Q(divisor_q[45]) );
  DFF_X1 divisor_q_reg_43_ ( .D(n532), .CK(clk_i), .Q(divisor_q[43]) );
  DFF_X1 divisor_q_reg_42_ ( .D(n533), .CK(clk_i), .Q(divisor_q[42]) );
  DFF_X1 divisor_q_reg_40_ ( .D(n535), .CK(clk_i), .Q(divisor_q[40]) );
  DFF_X1 divisor_q_reg_35_ ( .D(n540), .CK(clk_i), .Q(divisor_q[35]) );
  DFF_X1 divisor_q_reg_34_ ( .D(n541), .CK(clk_i), .Q(divisor_q[34]) );
  DFF_X1 divisor_q_reg_32_ ( .D(n543), .CK(clk_i), .Q(divisor_q[32]) );
  DFF_X1 divisor_q_reg_44_ ( .D(n531), .CK(clk_i), .Q(divisor_q[44]) );
  DFF_X1 divisor_q_reg_41_ ( .D(n534), .CK(clk_i), .Q(divisor_q[41]) );
  DFF_X1 divisor_q_reg_39_ ( .D(n536), .CK(clk_i), .Q(divisor_q[39]) );
  DFF_X1 divisor_q_reg_38_ ( .D(n537), .CK(clk_i), .Q(divisor_q[38]) );
  DFF_X1 divisor_q_reg_37_ ( .D(n538), .CK(clk_i), .Q(divisor_q[37]) );
  DFF_X1 divisor_q_reg_36_ ( .D(n539), .CK(clk_i), .Q(divisor_q[36]) );
  DFF_X1 divisor_q_reg_31_ ( .D(n544), .CK(clk_i), .Q(divisor_q[31]) );
  DFF_X1 divisor_q_reg_46_ ( .D(n529), .CK(clk_i), .Q(divisor_q[46]) );
  DFF_X1 divisor_q_reg_47_ ( .D(n528), .CK(clk_i), .Q(divisor_q[47]) );
  DFF_X1 divisor_q_reg_48_ ( .D(n527), .CK(clk_i), .Q(divisor_q[48]) );
  DFF_X1 divisor_q_reg_49_ ( .D(n526), .CK(clk_i), .Q(divisor_q[49]) );
  DFF_X1 divisor_q_reg_50_ ( .D(n525), .CK(clk_i), .Q(divisor_q[50]) );
  DFF_X1 divisor_q_reg_51_ ( .D(n524), .CK(clk_i), .Q(divisor_q[51]) );
  DFF_X1 divisor_q_reg_52_ ( .D(n523), .CK(clk_i), .Q(divisor_q[52]) );
  DFF_X1 divisor_q_reg_53_ ( .D(n522), .CK(clk_i), .Q(divisor_q[53]) );
  DFF_X1 divisor_q_reg_54_ ( .D(n521), .CK(clk_i), .Q(divisor_q[54]) );
  DFF_X1 divisor_q_reg_55_ ( .D(n520), .CK(clk_i), .Q(divisor_q[55]) );
  DFF_X1 divisor_q_reg_56_ ( .D(n519), .CK(clk_i), .Q(divisor_q[56]) );
  DFF_X1 divisor_q_reg_57_ ( .D(n518), .CK(clk_i), .Q(divisor_q[57]) );
  DFF_X1 divisor_q_reg_58_ ( .D(n517), .CK(clk_i), .Q(divisor_q[58]) );
  DFF_X1 divisor_q_reg_59_ ( .D(n516), .CK(clk_i), .Q(divisor_q[59]) );
  DFF_X1 divisor_q_reg_60_ ( .D(n515), .CK(clk_i), .Q(divisor_q[60]) );
  DFF_X1 divisor_q_reg_61_ ( .D(n514), .CK(clk_i), .Q(divisor_q[61]) );
  DFF_X1 result_q_reg_0_ ( .D(n417), .CK(clk_i), .Q(result_o[0]) );
  DFF_X1 result_q_reg_4_ ( .D(n421), .CK(clk_i), .Q(result_o[4]) );
  DFF_X1 result_q_reg_3_ ( .D(n420), .CK(clk_i), .Q(result_o[3]) );
  DFF_X1 result_q_reg_5_ ( .D(n422), .CK(clk_i), .Q(result_o[5]) );
  DFF_X1 result_q_reg_6_ ( .D(n423), .CK(clk_i), .Q(result_o[6]) );
  DFF_X1 result_q_reg_7_ ( .D(n424), .CK(clk_i), .Q(result_o[7]) );
  DFF_X1 result_q_reg_12_ ( .D(n429), .CK(clk_i), .Q(result_o[12]) );
  DFF_X1 result_q_reg_9_ ( .D(n426), .CK(clk_i), .Q(result_o[9]) );
  DFF_X1 result_q_reg_8_ ( .D(n425), .CK(clk_i), .Q(result_o[8]) );
  DFF_X1 result_q_reg_10_ ( .D(n427), .CK(clk_i), .Q(result_o[10]) );
  DFF_X1 result_q_reg_13_ ( .D(n430), .CK(clk_i), .Q(result_o[13]) );
  DFF_X1 result_q_reg_15_ ( .D(n432), .CK(clk_i), .Q(result_o[15]) );
  DFF_X1 result_q_reg_11_ ( .D(n428), .CK(clk_i), .Q(result_o[11]) );
  DFF_X1 result_q_reg_14_ ( .D(n431), .CK(clk_i), .Q(result_o[14]) );
  DFF_X1 result_q_reg_16_ ( .D(n433), .CK(clk_i), .Q(result_o[16]) );
  DFF_X1 result_q_reg_17_ ( .D(n434), .CK(clk_i), .Q(result_o[17]) );
  DFF_X1 result_q_reg_18_ ( .D(n435), .CK(clk_i), .Q(result_o[18]) );
  DFF_X1 result_q_reg_19_ ( .D(n436), .CK(clk_i), .Q(result_o[19]) );
  DFF_X1 result_q_reg_20_ ( .D(n437), .CK(clk_i), .Q(result_o[20]) );
  DFF_X1 result_q_reg_21_ ( .D(n438), .CK(clk_i), .Q(result_o[21]) );
  DFF_X1 result_q_reg_22_ ( .D(n439), .CK(clk_i), .Q(result_o[22]) );
  DFF_X1 result_q_reg_23_ ( .D(n440), .CK(clk_i), .Q(result_o[23]) );
  DFF_X1 result_q_reg_27_ ( .D(n444), .CK(clk_i), .Q(result_o[27]) );
  DFF_X1 result_q_reg_28_ ( .D(n445), .CK(clk_i), .Q(result_o[28]) );
  DFF_X1 result_q_reg_26_ ( .D(n443), .CK(clk_i), .Q(result_o[26]) );
  DFF_X1 result_q_reg_25_ ( .D(n442), .CK(clk_i), .Q(result_o[25]) );
  DFF_X1 result_q_reg_31_ ( .D(n448), .CK(clk_i), .Q(result_o[31]) );
  DFF_X1 result_q_reg_24_ ( .D(n441), .CK(clk_i), .Q(result_o[24]) );
  DFF_X2 mul_operand_b_q_reg_23_ ( .D(N79), .CK(clk_i), .Q(mul_operand_b_q[23]) );
  DFF_X2 mul_operand_b_q_reg_29_ ( .D(N85), .CK(clk_i), .Q(mul_operand_b_q[29]), .QN(n985) );
  DFF_X2 mul_operand_b_q_reg_27_ ( .D(N83), .CK(clk_i), .Q(mul_operand_b_q[27]), .QN(n837) );
  DFF_X2 mul_operand_b_q_reg_22_ ( .D(N78), .CK(clk_i), .Q(mul_operand_b_q[22]) );
  DFF_X2 mul_operand_b_q_reg_25_ ( .D(N81), .CK(clk_i), .Q(mul_operand_b_q[25]) );
  DFF_X2 mul_operand_b_q_reg_21_ ( .D(N77), .CK(clk_i), .Q(mul_operand_b_q[21]) );
  DFF_X2 mul_operand_b_q_reg_18_ ( .D(N74), .CK(clk_i), .Q(mul_operand_b_q[18]), .QN(n347) );
  DFF_X2 mul_operand_b_q_reg_12_ ( .D(N68), .CK(clk_i), .Q(mul_operand_b_q[12]), .QN(n349) );
  DFF_X2 mul_operand_b_q_reg_15_ ( .D(N71), .CK(clk_i), .Q(mul_operand_b_q[15]) );
  DFF_X2 mul_operand_a_q_reg_32_ ( .D(n402), .CK(clk_i), .QN(
        mul_operand_a_q[32]) );
  SDFF_X2 mul_operand_a_q_reg_23_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[23]), 
        .CK(clk_i), .Q(mul_operand_a_q[23]) );
  SDFF_X2 mul_operand_a_q_reg_26_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[26]), 
        .CK(clk_i), .Q(mul_operand_a_q[26]) );
  SDFF_X2 mul_operand_a_q_reg_29_ ( .D(1'b0), .SI(n611), .SE(operand_ra_i[29]), 
        .CK(clk_i), .Q(mul_operand_a_q[29]) );
  DFF_X2 mul_operand_b_q_reg_17_ ( .D(N73), .CK(clk_i), .Q(mul_operand_b_q[17]), .QN(n350) );
  DFF_X2 mul_operand_b_q_reg_13_ ( .D(N69), .CK(clk_i), .Q(mul_operand_b_q[13]) );
  DFF_X2 mul_operand_b_q_reg_7_ ( .D(N63), .CK(clk_i), .Q(mul_operand_b_q[7])
         );
  DFF_X2 mul_operand_b_q_reg_20_ ( .D(N76), .CK(clk_i), .Q(mul_operand_b_q[20]), .QN(n2369) );
  DFF_X2 mul_operand_b_q_reg_11_ ( .D(N67), .CK(clk_i), .Q(mul_operand_b_q[11]) );
  DFF_X2 mul_operand_b_q_reg_4_ ( .D(N60), .CK(clk_i), .Q(mul_operand_b_q[4])
         );
  DFF_X2 mul_operand_b_q_reg_8_ ( .D(N64), .CK(clk_i), .Q(mul_operand_b_q[8])
         );
  DFF_X2 mul_operand_b_q_reg_14_ ( .D(N70), .CK(clk_i), .Q(mul_operand_b_q[14]) );
  DFF_X2 mul_operand_b_q_reg_10_ ( .D(N66), .CK(clk_i), .Q(mul_operand_b_q[10]) );
  DFF_X2 mul_operand_b_q_reg_19_ ( .D(N75), .CK(clk_i), .Q(mul_operand_b_q[19]), .QN(n2366) );
  AOI21_X1 U3 ( .B1(mult_x_6_n278), .B2(n932), .A(n877), .ZN(n931) );
  INV_X1 U4 ( .A(n941), .ZN(mult_x_6_n286) );
  AND2_X1 U5 ( .A1(n1963), .A2(n2049), .ZN(n2047) );
  XOR2_X1 U6 ( .A(mult_x_6_n1063), .B(n2247), .Z(mult_x_6_n1095) );
  BUF_X1 U7 ( .A(mul_operand_a_q[5]), .Z(n2176) );
  BUF_X2 U8 ( .A(mul_operand_b_q[4]), .Z(n2192) );
  INV_X1 U9 ( .A(n2178), .ZN(n2179) );
  INV_X1 U10 ( .A(n931), .ZN(mult_x_6_n277) );
  XNOR2_X1 U11 ( .A(mult_x_6_n278), .B(n930), .ZN(mult_result_w[53]) );
  XNOR2_X1 U12 ( .A(mult_x_6_n857), .B(mult_x_6_n1462), .ZN(n804) );
  XNOR2_X1 U13 ( .A(mult_x_6_n312), .B(n928), .ZN(mult_result_w[19]) );
  INV_X1 U14 ( .A(n933), .ZN(mult_x_6_n280) );
  XNOR2_X1 U15 ( .A(mult_x_6_n283), .B(n898), .ZN(mult_result_w[48]) );
  XNOR2_X1 U16 ( .A(mult_x_6_n945), .B(mult_x_6_n1470), .ZN(n861) );
  AOI222_X1 U17 ( .A1(mult_x_6_n1103), .A2(n1665), .B1(n2195), .B2(n1666), 
        .C1(n1018), .C2(n2203), .ZN(n1) );
  XOR2_X1 U18 ( .A(n2171), .B(n1), .Z(n2) );
  INV_X1 U19 ( .A(mult_x_6_n934), .ZN(n3) );
  NOR2_X1 U20 ( .A1(n2), .A2(n3), .ZN(mult_x_6_n924) );
  XNOR2_X1 U21 ( .A(n2), .B(mult_x_6_n934), .ZN(mult_x_6_n925) );
  INV_X1 U22 ( .A(n2171), .ZN(n4) );
  AOI21_X1 U23 ( .B1(n2149), .B2(n2196), .A(n4), .ZN(mult_x_6_n934) );
  AND2_X1 U24 ( .A1(n2149), .A2(n2196), .ZN(mult_x_6_n935) );
  AOI22_X1 U25 ( .A1(mult_x_6_n1102), .A2(n2214), .B1(n2145), .B2(n2196), .ZN(
        n5) );
  AOI22_X1 U26 ( .A1(n1959), .A2(n1009), .B1(n2195), .B2(n2216), .ZN(n6) );
  NAND2_X1 U27 ( .A1(n6), .A2(n5), .ZN(n7) );
  XNOR2_X1 U28 ( .A(n7), .B(n348), .ZN(mult_x_6_n1411) );
  AND3_X2 U29 ( .A1(n2143), .A2(n19601), .A3(n1963), .ZN(n2144) );
  AOI222_X1 U30 ( .A1(n1958), .A2(mult_x_6_n1103), .B1(n2196), .B2(n2216), 
        .C1(n2286), .C2(n1959), .ZN(n8) );
  XNOR2_X1 U31 ( .A(n8), .B(n348), .ZN(n9) );
  INV_X1 U32 ( .A(mult_x_6_n988), .ZN(n10) );
  NOR2_X1 U33 ( .A1(n9), .A2(n10), .ZN(mult_x_6_n984) );
  XNOR2_X1 U34 ( .A(mult_x_6_n988), .B(n9), .ZN(mult_x_6_n985) );
  AND2_X1 U35 ( .A1(n985), .A2(n353), .ZN(n11) );
  OR2_X1 U36 ( .A1(n983), .A2(n11), .ZN(n12) );
  OAI222_X1 U37 ( .A1(n12), .A2(n984), .B1(n985), .B2(n353), .C1(n11), .C2(
        n2275), .ZN(mult_x_6_n1042) );
  INV_X1 U38 ( .A(mult_x_6_n1425), .ZN(n13) );
  INV_X1 U39 ( .A(mult_x_6_n783), .ZN(n14) );
  OAI21_X1 U40 ( .B1(mult_x_6_n783), .B2(mult_x_6_n1425), .A(n801), .ZN(n15)
         );
  OAI21_X1 U41 ( .B1(n13), .B2(n14), .A(n15), .ZN(n693) );
  NAND3_X1 U42 ( .A1(n2259), .A2(n2257), .A3(n2258), .ZN(n16) );
  OAI222_X1 U43 ( .A1(n16), .A2(n2194), .B1(n16), .B2(mul_operand_b_q[4]), 
        .C1(n2194), .C2(mul_operand_b_q[4]), .ZN(n17) );
  INV_X1 U44 ( .A(n17), .ZN(mult_x_6_n1067) );
  AOI222_X1 U45 ( .A1(n2196), .A2(n2205), .B1(n1767), .B2(mult_x_6_n1103), 
        .C1(n2195), .C2(n2208), .ZN(n18) );
  XOR2_X1 U46 ( .A(n2172), .B(n18), .Z(n19) );
  INV_X1 U47 ( .A(mult_x_6_n958), .ZN(n20) );
  NOR2_X1 U48 ( .A1(n19), .A2(n20), .ZN(mult_x_6_n950) );
  XNOR2_X1 U49 ( .A(n19), .B(mult_x_6_n958), .ZN(mult_x_6_n951) );
  INV_X1 U50 ( .A(mul_operand_b_q[29]), .ZN(n21) );
  INV_X1 U51 ( .A(mult_x_6_n1042), .ZN(n22) );
  OAI21_X1 U52 ( .B1(mul_operand_b_q[29]), .B2(mult_x_6_n1042), .A(
        mul_operand_b_q[30]), .ZN(n23) );
  OAI21_X1 U53 ( .B1(n21), .B2(n22), .A(n23), .ZN(mult_x_6_n1041) );
  INV_X1 U54 ( .A(mult_x_6_n1430), .ZN(n24) );
  INV_X1 U55 ( .A(mult_x_6_n859), .ZN(n25) );
  OAI21_X1 U56 ( .B1(mult_x_6_n859), .B2(mult_x_6_n1430), .A(mult_x_6_n870), 
        .ZN(n26) );
  OAI21_X1 U57 ( .B1(n24), .B2(n25), .A(n26), .ZN(mult_x_6_n856) );
  OAI21_X1 U58 ( .B1(mult_x_6_n947), .B2(n2359), .A(n757), .ZN(n2360) );
  AOI222_X1 U59 ( .A1(n2142), .A2(n2193), .B1(n1009), .B2(n608), .C1(n2286), 
        .C2(n2119), .ZN(n27) );
  NAND2_X1 U60 ( .A1(n2120), .A2(mult_x_6_n1101), .ZN(n28) );
  NAND2_X1 U61 ( .A1(n28), .A2(n27), .ZN(n29) );
  XNOR2_X1 U62 ( .A(n29), .B(n1013), .ZN(mult_x_6_n1480) );
  INV_X1 U63 ( .A(mult_x_6_n1330), .ZN(n30) );
  INV_X1 U64 ( .A(mult_x_6_n805), .ZN(n31) );
  OAI21_X1 U65 ( .B1(mult_x_6_n805), .B2(mult_x_6_n1330), .A(n698), .ZN(n32)
         );
  OAI21_X1 U66 ( .B1(n30), .B2(n31), .A(n32), .ZN(mult_x_6_n802) );
  INV_X1 U67 ( .A(mult_x_6_n1374), .ZN(n33) );
  INV_X1 U68 ( .A(mult_x_6_n951), .ZN(n34) );
  OAI21_X1 U69 ( .B1(mult_x_6_n951), .B2(mult_x_6_n1374), .A(mult_x_6_n956), 
        .ZN(n35) );
  OAI21_X1 U70 ( .B1(n33), .B2(n34), .A(n35), .ZN(mult_x_6_n948) );
  AOI222_X1 U71 ( .A1(n2190), .A2(n2218), .B1(n2192), .B2(n1020), .C1(n2193), 
        .C2(n2145), .ZN(n36) );
  NAND2_X1 U72 ( .A1(n2214), .A2(n355), .ZN(n37) );
  NAND2_X1 U73 ( .A1(n36), .A2(n37), .ZN(n38) );
  XOR2_X1 U74 ( .A(n2174), .B(n38), .Z(mult_x_6_n1408) );
  INV_X1 U75 ( .A(n949), .ZN(n39) );
  NOR2_X1 U76 ( .A1(n6701), .A2(n39), .ZN(n667) );
  AOI22_X1 U77 ( .A1(mult_x_6_n333), .A2(mult_x_6_n334), .B1(n2305), .B2(n2307), .ZN(n40) );
  OAI21_X1 U78 ( .B1(n2240), .B2(n2304), .A(n40), .ZN(n2428) );
  XNOR2_X1 U79 ( .A(mult_x_6_n1425), .B(n801), .ZN(n41) );
  XNOR2_X1 U80 ( .A(n41), .B(mult_x_6_n783), .ZN(mult_x_6_n781) );
  AND2_X1 U81 ( .A1(n2049), .A2(n2196), .ZN(mult_x_6_n995) );
  INV_X1 U82 ( .A(n2176), .ZN(n42) );
  AOI21_X1 U83 ( .B1(n2049), .B2(n2196), .A(n42), .ZN(mult_x_6_n994) );
  AOI222_X1 U84 ( .A1(mult_x_6_n803), .A2(mult_x_6_n816), .B1(mult_x_6_n803), 
        .B2(mult_x_6_n1362), .C1(mult_x_6_n816), .C2(mult_x_6_n1362), .ZN(n847) );
  AOI22_X1 U85 ( .A1(n1020), .A2(n2193), .B1(n2217), .B2(mul_operand_b_q[4]), 
        .ZN(n43) );
  AOI22_X1 U86 ( .A1(n1009), .A2(n405), .B1(n2214), .B2(n622), .ZN(n44) );
  NAND2_X1 U87 ( .A1(n44), .A2(n43), .ZN(n45) );
  XNOR2_X1 U88 ( .A(n45), .B(n348), .ZN(mult_x_6_n1409) );
  AOI22_X1 U89 ( .A1(mult_x_6_n340), .A2(mult_x_6_n337), .B1(n950), .B2(n951), 
        .ZN(n46) );
  INV_X1 U90 ( .A(n46), .ZN(n948) );
  NOR2_X1 U91 ( .A1(mult_x_6_n1437), .A2(mult_x_6_n939), .ZN(n47) );
  NAND2_X1 U92 ( .A1(mult_x_6_n1437), .A2(mult_x_6_n939), .ZN(n48) );
  OAI221_X1 U93 ( .B1(n47), .B2(n2355), .C1(n47), .C2(n2360), .A(n48), .ZN(
        mult_x_6_n936) );
  AOI222_X1 U94 ( .A1(n2223), .A2(n2190), .B1(n2221), .B2(n2192), .C1(n2193), 
        .C2(n2144), .ZN(n49) );
  NAND2_X1 U95 ( .A1(n2219), .A2(n1024), .ZN(n50) );
  NAND2_X1 U96 ( .A1(n50), .A2(n49), .ZN(n51) );
  XNOR2_X1 U97 ( .A(n51), .B(n1026), .ZN(mult_x_6_n1443) );
  NOR2_X1 U98 ( .A1(n935), .A2(n2408), .ZN(n52) );
  AOI21_X1 U99 ( .B1(mult_x_6_n520), .B2(mult_x_6_n506), .A(n52), .ZN(n644) );
  OAI21_X1 U100 ( .B1(mult_x_6_n1419), .B2(mult_x_6_n669), .A(mult_x_6_n686), 
        .ZN(n2345) );
  AOI222_X1 U101 ( .A1(n2195), .A2(n2141), .B1(n1009), .B2(n2142), .C1(n2196), 
        .C2(n2119), .ZN(n53) );
  NAND2_X1 U102 ( .A1(n2120), .A2(mult_x_6_n1102), .ZN(n54) );
  NAND2_X1 U103 ( .A1(n54), .A2(n53), .ZN(n55) );
  XNOR2_X1 U104 ( .A(n55), .B(n1013), .ZN(mult_x_6_n1481) );
  AOI22_X1 U105 ( .A1(n2581), .A2(dividend_q[26]), .B1(n2580), .B2(
        result_o[26]), .ZN(n5610) );
  XOR2_X1 U106 ( .A(mult_x_6_n346), .B(mult_x_6_n344), .Z(n579) );
  OAI21_X1 U107 ( .B1(mult_x_6_n273), .B2(n579), .A(n2993), .ZN(n581) );
  AOI21_X1 U108 ( .B1(mult_x_6_n273), .B2(n579), .A(n581), .ZN(n590) );
  XOR2_X1 U109 ( .A(mult_x_6_n781), .B(mult_x_6_n1457), .Z(n600) );
  OAI21_X1 U110 ( .B1(n8001), .B2(n600), .A(n2579), .ZN(n6100) );
  AOI21_X1 U111 ( .B1(n8001), .B2(n600), .A(n6100), .ZN(n620) );
  AOI211_X1 U112 ( .C1(n2571), .C2(C22_DATA3_26), .A(n590), .B(n620), .ZN(
        n6300) );
  OAI211_X1 U113 ( .C1(n2799), .C2(n7700), .A(n5610), .B(n6300), .ZN(n443) );
  INV_X1 U114 ( .A(n2172), .ZN(n6500) );
  AOI21_X1 U115 ( .B1(n2147), .B2(n2196), .A(n6500), .ZN(mult_x_6_n958) );
  AND2_X1 U116 ( .A1(n2147), .A2(n2196), .ZN(mult_x_6_n959) );
  AOI222_X1 U117 ( .A1(n1009), .A2(n2144), .B1(n2221), .B2(n2193), .C1(n2222), 
        .C2(mul_operand_b_q[4]), .ZN(n695) );
  INV_X1 U118 ( .A(mult_x_6_n963), .ZN(n6600) );
  INV_X1 U119 ( .A(mult_x_6_n1440), .ZN(n6700) );
  OAI21_X1 U120 ( .B1(mult_x_6_n963), .B2(mult_x_6_n1440), .A(mult_x_6_n966), 
        .ZN(n6800) );
  OAI21_X1 U121 ( .B1(n6600), .B2(n6700), .A(n6800), .ZN(mult_x_6_n960) );
  INV_X1 U122 ( .A(n2307), .ZN(n6900) );
  OAI21_X1 U123 ( .B1(n2310), .B2(n2304), .A(n6900), .ZN(n2415) );
  OAI21_X1 U124 ( .B1(mult_x_6_n341), .B2(n2302), .A(n2254), .ZN(n7000) );
  OAI21_X1 U125 ( .B1(n105), .B2(n106), .A(n7000), .ZN(n951) );
  INV_X1 U126 ( .A(mult_x_6_n343), .ZN(n105) );
  INV_X1 U127 ( .A(mult_x_6_n341), .ZN(n106) );
  XNOR2_X1 U128 ( .A(n693), .B(mult_x_6_n765), .ZN(n107) );
  XNOR2_X1 U129 ( .A(n107), .B(mult_x_6_n1424), .ZN(mult_x_6_n763) );
  OR2_X1 U130 ( .A1(n2142), .A2(n2141), .ZN(n108) );
  AOI222_X1 U131 ( .A1(n108), .A2(mul_operand_b_q[32]), .B1(n2225), .B2(
        mult_x_6_n1071), .C1(n2179), .C2(n2224), .ZN(n109) );
  XNOR2_X1 U132 ( .A(mul_operand_a_q[2]), .B(n109), .ZN(mult_x_6_n1450) );
  NAND2_X1 U133 ( .A1(result_o[18]), .A2(n2580), .ZN(n110) );
  OAI21_X1 U134 ( .B1(n8500), .B2(n2799), .A(n110), .ZN(n111) );
  AOI21_X1 U135 ( .B1(dividend_q[18]), .B2(n2581), .A(n111), .ZN(n112) );
  AOI22_X1 U136 ( .A1(C22_DATA3_18), .A2(n2571), .B1(n2579), .B2(
        mult_result_w[18]), .ZN(n113) );
  XOR2_X1 U137 ( .A(mult_x_6_n281), .B(mult_x_6_n404), .Z(n114) );
  NAND2_X1 U138 ( .A1(mult_x_6_n396), .A2(n114), .ZN(n115) );
  OAI211_X1 U139 ( .C1(mult_x_6_n396), .C2(n114), .A(n115), .B(n2578), .ZN(
        n116) );
  NAND3_X1 U140 ( .A1(n112), .A2(n113), .A3(n116), .ZN(n435) );
  AOI22_X1 U141 ( .A1(n2581), .A2(dividend_q[9]), .B1(n2580), .B2(result_o[9]), 
        .ZN(n117) );
  XOR2_X1 U142 ( .A(mult_x_6_n506), .B(mult_x_6_n520), .Z(n118) );
  OAI21_X1 U143 ( .B1(n2339), .B2(n2338), .A(n2408), .ZN(n119) );
  OAI21_X1 U144 ( .B1(n118), .B2(n119), .A(n2578), .ZN(n120) );
  AOI21_X1 U145 ( .B1(n118), .B2(n119), .A(n120), .ZN(n121) );
  XOR2_X1 U146 ( .A(mult_x_6_n1474), .B(mult_x_6_n973), .Z(n122) );
  OAI21_X1 U147 ( .B1(n753), .B2(n122), .A(n2579), .ZN(n123) );
  AOI21_X1 U148 ( .B1(n753), .B2(n122), .A(n123), .ZN(n124) );
  AOI211_X1 U149 ( .C1(n2800), .C2(C22_DATA3_9), .A(n121), .B(n124), .ZN(n125)
         );
  OAI211_X1 U150 ( .C1(n2799), .C2(n94), .A(n117), .B(n125), .ZN(n426) );
  NAND2_X1 U151 ( .A1(n2581), .A2(dividend_q[5]), .ZN(n126) );
  OAI21_X1 U152 ( .B1(n98), .B2(n2799), .A(n126), .ZN(n127) );
  AOI21_X1 U153 ( .B1(result_o[5]), .B2(n2580), .A(n127), .ZN(n128) );
  AOI22_X1 U154 ( .A1(C22_DATA3_5), .A2(n2571), .B1(n2994), .B2(
        mult_result_w[5]), .ZN(n129) );
  XOR2_X1 U155 ( .A(mult_x_6_n294), .B(mult_x_6_n588), .Z(n130) );
  NAND2_X1 U156 ( .A1(mult_x_6_n571), .A2(n130), .ZN(n131) );
  OAI211_X1 U157 ( .C1(mult_x_6_n571), .C2(n130), .A(n131), .B(n2578), .ZN(
        n132) );
  NAND3_X1 U158 ( .A1(n128), .A2(n129), .A3(n132), .ZN(n422) );
  AOI222_X1 U159 ( .A1(mult_x_6_n849), .A2(mult_x_6_n860), .B1(mult_x_6_n849), 
        .B2(mult_x_6_n1365), .C1(mult_x_6_n860), .C2(mult_x_6_n1365), .ZN(n818) );
  AOI222_X1 U160 ( .A1(mult_x_6_n789), .A2(mult_x_6_n802), .B1(mult_x_6_n789), 
        .B2(mult_x_6_n1329), .C1(mult_x_6_n802), .C2(mult_x_6_n1329), .ZN(n772) );
  AOI222_X1 U161 ( .A1(n2196), .A2(n2211), .B1(n1868), .B2(mult_x_6_n1103), 
        .C1(n2195), .C2(n2212), .ZN(n133) );
  XNOR2_X1 U162 ( .A(n133), .B(n633), .ZN(n134) );
  INV_X1 U163 ( .A(mult_x_6_n976), .ZN(n135) );
  NOR2_X1 U164 ( .A1(n134), .A2(n135), .ZN(mult_x_6_n970) );
  XNOR2_X1 U165 ( .A(mult_x_6_n976), .B(n134), .ZN(mult_x_6_n971) );
  AOI222_X1 U166 ( .A1(n2221), .A2(n2190), .B1(n2144), .B2(mul_operand_b_q[4]), 
        .C1(n2222), .C2(n2189), .ZN(n136) );
  INV_X1 U167 ( .A(n136), .ZN(n857) );
  XNOR2_X1 U168 ( .A(mult_x_6_n1431), .B(mult_x_6_n882), .ZN(n137) );
  XNOR2_X1 U169 ( .A(n137), .B(mult_x_6_n873), .ZN(mult_x_6_n871) );
  XNOR2_X1 U170 ( .A(mult_x_6_n1435), .B(mult_x_6_n926), .ZN(n138) );
  XNOR2_X1 U171 ( .A(n138), .B(mult_x_6_n919), .ZN(mult_x_6_n917) );
  AOI22_X1 U172 ( .A1(n2581), .A2(dividend_q[30]), .B1(n2580), .B2(
        result_o[30]), .ZN(n139) );
  OAI21_X1 U173 ( .B1(n2799), .B2(n7300), .A(n139), .ZN(n140) );
  AOI21_X1 U174 ( .B1(n2571), .B2(C22_DATA3_30), .A(n140), .ZN(n141) );
  XOR2_X1 U175 ( .A(mult_x_6_n301), .B(mult_x_6_n1453), .Z(n142) );
  NAND2_X1 U176 ( .A1(mult_x_6_n707), .A2(n142), .ZN(n143) );
  OAI211_X1 U177 ( .C1(mult_x_6_n707), .C2(n142), .A(n2579), .B(n143), .ZN(
        n144) );
  NAND2_X1 U178 ( .A1(n141), .A2(n144), .ZN(n609) );
  INV_X1 U179 ( .A(mult_x_6_n270), .ZN(n145) );
  NAND3_X1 U180 ( .A1(n2578), .A2(n946), .A3(n145), .ZN(n146) );
  INV_X1 U181 ( .A(n387), .ZN(n147) );
  NAND4_X1 U182 ( .A1(n1001), .A2(mult_x_6_n270), .A3(n2415), .A4(n147), .ZN(
        n148) );
  OR2_X1 U183 ( .A1(n997), .A2(n999), .ZN(n149) );
  NAND4_X1 U184 ( .A1(n2528), .A2(n146), .A3(n148), .A4(n149), .ZN(n448) );
  AOI22_X1 U185 ( .A1(n2580), .A2(result_o[8]), .B1(dividend_q[8]), .B2(n2581), 
        .ZN(n150) );
  XNOR2_X1 U186 ( .A(mult_x_6_n535), .B(mult_x_6_n521), .ZN(n151) );
  OAI21_X1 U187 ( .B1(n2339), .B2(n151), .A(n2578), .ZN(n152) );
  AOI21_X1 U188 ( .B1(n2339), .B2(n151), .A(n152), .ZN(n153) );
  XOR2_X1 U189 ( .A(mult_x_6_n1475), .B(mult_x_6_n979), .Z(n154) );
  OAI21_X1 U190 ( .B1(mult_x_6_n323), .B2(n154), .A(n2579), .ZN(n155) );
  AOI21_X1 U191 ( .B1(mult_x_6_n323), .B2(n154), .A(n155), .ZN(n156) );
  AOI211_X1 U192 ( .C1(n2800), .C2(C22_DATA3_8), .A(n153), .B(n156), .ZN(n157)
         );
  OAI211_X1 U193 ( .C1(n2799), .C2(n95), .A(n150), .B(n157), .ZN(n425) );
  INV_X1 U194 ( .A(mul_operand_b_q[23]), .ZN(n158) );
  INV_X1 U195 ( .A(mult_x_6_n1049), .ZN(n159) );
  OAI21_X1 U196 ( .B1(mul_operand_b_q[23]), .B2(mult_x_6_n1049), .A(
        mul_operand_b_q[22]), .ZN(n160) );
  OAI21_X1 U197 ( .B1(n158), .B2(n159), .A(n160), .ZN(n2250) );
  XOR2_X1 U198 ( .A(mult_x_6_n1358), .B(mult_x_6_n733), .Z(n161) );
  XNOR2_X1 U199 ( .A(n8501), .B(n161), .ZN(mult_x_6_n731) );
  XOR2_X1 U200 ( .A(mult_x_6_n1067), .B(n2285), .Z(n1024) );
  INV_X1 U201 ( .A(n2412), .ZN(n162) );
  AOI22_X1 U202 ( .A1(mult_x_6_n352), .A2(mult_x_6_n347), .B1(n917), .B2(n162), 
        .ZN(n6701) );
  NAND3_X1 U203 ( .A1(n2245), .A2(n2322), .A3(n2246), .ZN(n163) );
  NAND2_X1 U204 ( .A1(n163), .A2(n2321), .ZN(n164) );
  XOR2_X1 U205 ( .A(mul_operand_b_q[10]), .B(mul_operand_b_q[11]), .Z(n165) );
  XNOR2_X1 U206 ( .A(n164), .B(n165), .ZN(mult_x_6_n1093) );
  OAI21_X1 U207 ( .B1(mult_x_6_n960), .B2(mult_x_6_n955), .A(mult_x_6_n1439), 
        .ZN(n166) );
  OAI21_X1 U208 ( .B1(n167), .B2(n168), .A(n166), .ZN(n757) );
  INV_X1 U209 ( .A(mult_x_6_n960), .ZN(n167) );
  INV_X1 U210 ( .A(mult_x_6_n955), .ZN(n168) );
  NOR2_X1 U211 ( .A1(mult_x_6_n476), .A2(mult_x_6_n489), .ZN(n169) );
  AOI21_X1 U212 ( .B1(n2343), .B2(n2413), .A(n169), .ZN(n1005) );
  AOI22_X1 U213 ( .A1(mult_x_6_n1102), .A2(n2047), .B1(n2144), .B2(n2196), 
        .ZN(n17000) );
  OAI211_X1 U214 ( .C1(n2046), .C2(n963), .A(n958), .B(n959), .ZN(n17100) );
  AOI21_X1 U215 ( .B1(n962), .B2(n17000), .A(n17100), .ZN(n17200) );
  INV_X1 U216 ( .A(n17200), .ZN(n964) );
  AOI222_X1 U217 ( .A1(mult_x_6_n671), .A2(mult_x_6_n688), .B1(mult_x_6_n671), 
        .B2(mult_x_6_n1387), .C1(mult_x_6_n688), .C2(mult_x_6_n1387), .ZN(
        n2379) );
  XNOR2_X1 U218 ( .A(mult_x_6_n969), .B(mult_x_6_n972), .ZN(n17300) );
  XNOR2_X1 U219 ( .A(n17300), .B(mult_x_6_n1441), .ZN(mult_x_6_n967) );
  XNOR2_X1 U220 ( .A(mult_x_6_n337), .B(mult_x_6_n340), .ZN(n17400) );
  AOI21_X1 U221 ( .B1(mult_x_6_n273), .B2(n2303), .A(n951), .ZN(n17500) );
  XNOR2_X1 U222 ( .A(n17500), .B(n17400), .ZN(n17600) );
  OAI21_X1 U223 ( .B1(n2799), .B2(n7500), .A(n2796), .ZN(n17700) );
  AOI21_X1 U224 ( .B1(n2571), .B2(C22_DATA3_28), .A(n17700), .ZN(n17800) );
  XOR2_X1 U225 ( .A(n881), .B(mult_x_6_n1455), .Z(n17900) );
  NAND2_X1 U226 ( .A1(mult_x_6_n745), .A2(n17900), .ZN(n18000) );
  OAI211_X1 U227 ( .C1(mult_x_6_n745), .C2(n17900), .A(n2579), .B(n18000), 
        .ZN(n18100) );
  OAI211_X1 U228 ( .C1(n17600), .C2(n387), .A(n17800), .B(n18100), .ZN(n445)
         );
  AOI22_X1 U229 ( .A1(dividend_q[0]), .A2(n2581), .B1(n2580), .B2(result_o[0]), 
        .ZN(n18200) );
  XNOR2_X1 U230 ( .A(mult_x_6_n1451), .B(mult_x_6_n299), .ZN(n18300) );
  XNOR2_X1 U231 ( .A(n18300), .B(mult_x_6_n667), .ZN(n18400) );
  AOI22_X1 U232 ( .A1(n2578), .A2(n18400), .B1(mult_result_w[0]), .B2(n2994), 
        .ZN(n18500) );
  INV_X1 U233 ( .A(n2799), .ZN(n18600) );
  INV_X1 U234 ( .A(n2746), .ZN(n18700) );
  AOI22_X1 U235 ( .A1(quotient_q[0]), .A2(n18600), .B1(n2571), .B2(n18700), 
        .ZN(n18800) );
  NAND3_X1 U236 ( .A1(n18200), .A2(n18500), .A3(n18800), .ZN(n417) );
  NOR4_X1 U237 ( .A1(operand_rb_i[11]), .A2(operand_rb_i[10]), .A3(
        operand_rb_i[9]), .A4(operand_rb_i[8]), .ZN(n18900) );
  NOR4_X1 U238 ( .A1(operand_rb_i[15]), .A2(operand_rb_i[14]), .A3(
        operand_rb_i[13]), .A4(operand_rb_i[12]), .ZN(n19000) );
  NOR4_X1 U239 ( .A1(operand_rb_i[3]), .A2(operand_rb_i[2]), .A3(
        operand_rb_i[1]), .A4(operand_rb_i[0]), .ZN(n19100) );
  NOR4_X1 U240 ( .A1(operand_rb_i[7]), .A2(operand_rb_i[6]), .A3(
        operand_rb_i[5]), .A4(operand_rb_i[4]), .ZN(n19200) );
  NAND4_X1 U241 ( .A1(n18900), .A2(n19000), .A3(n19100), .A4(n19200), .ZN(
        n19300) );
  NOR4_X1 U242 ( .A1(operand_rb_i[27]), .A2(operand_rb_i[26]), .A3(
        operand_rb_i[25]), .A4(operand_rb_i[24]), .ZN(n19400) );
  NOR4_X1 U243 ( .A1(operand_rb_i[31]), .A2(operand_rb_i[30]), .A3(
        operand_rb_i[29]), .A4(operand_rb_i[28]), .ZN(n19500) );
  NOR4_X1 U244 ( .A1(operand_rb_i[19]), .A2(operand_rb_i[18]), .A3(
        operand_rb_i[17]), .A4(operand_rb_i[16]), .ZN(n19600) );
  NOR4_X1 U245 ( .A1(operand_rb_i[23]), .A2(operand_rb_i[22]), .A3(
        operand_rb_i[21]), .A4(operand_rb_i[20]), .ZN(n19700) );
  NAND4_X1 U246 ( .A1(n19400), .A2(n19500), .A3(n19600), .A4(n19700), .ZN(
        n19800) );
  OAI22_X1 U247 ( .A1(n19300), .A2(n19800), .B1(operand_rb_i[31]), .B2(
        operand_ra_i[31]), .ZN(n19900) );
  AOI21_X1 U248 ( .B1(operand_rb_i[31]), .B2(operand_ra_i[31]), .A(n19900), 
        .ZN(n20000) );
  AOI22_X1 U249 ( .A1(operand_ra_i[31]), .A2(inst_rem_i), .B1(inst_div_i), 
        .B2(n20000), .ZN(n201) );
  OAI22_X1 U250 ( .A1(n2803), .A2(n201), .B1(n104), .B2(n2971), .ZN(n577) );
  INV_X1 U251 ( .A(mult_x_6_n1398), .ZN(n202) );
  INV_X1 U252 ( .A(mult_x_6_n861), .ZN(n203) );
  OAI21_X1 U253 ( .B1(mult_x_6_n861), .B2(mult_x_6_n1398), .A(mult_x_6_n872), 
        .ZN(n204) );
  OAI21_X1 U254 ( .B1(n202), .B2(n203), .A(n204), .ZN(mult_x_6_n858) );
  OAI21_X1 U255 ( .B1(mul_operand_b_q[17]), .B2(mult_x_6_n1055), .A(n2185), 
        .ZN(n205) );
  OAI21_X1 U256 ( .B1(n206), .B2(n207), .A(n205), .ZN(mult_x_6_n1054) );
  INV_X1 U257 ( .A(mul_operand_b_q[17]), .ZN(n206) );
  INV_X1 U258 ( .A(mult_x_6_n1055), .ZN(n207) );
  AOI222_X1 U259 ( .A1(n1020), .A2(n2190), .B1(n2226), .B2(mul_operand_b_q[4]), 
        .C1(n2217), .C2(n2188), .ZN(n208) );
  INV_X1 U260 ( .A(n208), .ZN(n817) );
  NAND3_X1 U261 ( .A1(n2284), .A2(n2392), .A3(n2283), .ZN(n209) );
  NAND2_X1 U262 ( .A1(n209), .A2(n2391), .ZN(n210) );
  XOR2_X1 U263 ( .A(n2189), .B(mul_operand_b_q[7]), .Z(n211) );
  XNOR2_X1 U264 ( .A(n210), .B(n211), .ZN(mult_x_6_n1097) );
  AOI22_X1 U265 ( .A1(n2179), .A2(n2132), .B1(mult_x_6_n1071), .B2(n2134), 
        .ZN(n212) );
  OAI21_X1 U266 ( .B1(n604), .B2(n632), .A(mul_operand_b_q[32]), .ZN(n213) );
  NAND2_X1 U267 ( .A1(n213), .A2(n212), .ZN(n214) );
  XNOR2_X1 U268 ( .A(n2122), .B(n214), .ZN(n2308) );
  OAI21_X1 U269 ( .B1(n2430), .B2(mult_x_6_n438), .A(mult_x_6_n448), .ZN(n215)
         );
  INV_X1 U270 ( .A(n215), .ZN(n2292) );
  XNOR2_X1 U271 ( .A(n2187), .B(mul_operand_b_q[10]), .ZN(n216) );
  NAND3_X1 U272 ( .A1(n2246), .A2(n2244), .A3(n2245), .ZN(n217) );
  XNOR2_X1 U273 ( .A(n217), .B(n216), .ZN(mult_x_6_n1094) );
  AOI222_X1 U274 ( .A1(mult_x_6_n1103), .A2(n2047), .B1(n2220), .B2(n2196), 
        .C1(n2048), .C2(n2286), .ZN(n218) );
  XOR2_X1 U275 ( .A(n218), .B(n1026), .Z(mult_x_6_n1447) );
  AOI22_X1 U276 ( .A1(dividend_q[31]), .A2(n2581), .B1(n2580), .B2(
        result_o[31]), .ZN(n219) );
  AOI22_X1 U277 ( .A1(dividend_q[31]), .A2(n2569), .B1(quotient_q[31]), .B2(
        n2570), .ZN(n220) );
  NAND2_X1 U278 ( .A1(DP_OP_63J3_127_9516_n1), .A2(n220), .ZN(n221) );
  OAI211_X1 U279 ( .C1(DP_OP_63J3_127_9516_n1), .C2(n220), .A(n221), .B(n2571), 
        .ZN(n222) );
  OAI211_X1 U280 ( .C1(n2799), .C2(n7200), .A(n219), .B(n222), .ZN(n223) );
  AOI21_X1 U281 ( .B1(n2579), .B2(mult_result_w[31]), .A(n223), .ZN(n2528) );
  XNOR2_X1 U282 ( .A(mult_x_6_n1436), .B(mult_x_6_n936), .ZN(n224) );
  XNOR2_X1 U283 ( .A(n224), .B(mult_x_6_n929), .ZN(mult_x_6_n927) );
  INV_X1 U284 ( .A(n1002), .ZN(n225) );
  INV_X1 U285 ( .A(n644), .ZN(n226) );
  AOI222_X1 U286 ( .A1(n225), .A2(n226), .B1(mult_x_6_n476), .B2(mult_x_6_n489), .C1(n1005), .C2(n1006), .ZN(n642) );
  INV_X1 U287 ( .A(mult_x_6_n1383), .ZN(n227) );
  INV_X1 U288 ( .A(mult_x_6_n1415), .ZN(n228) );
  OAI21_X1 U289 ( .B1(mult_x_6_n1415), .B2(mult_x_6_n1383), .A(mult_x_6_n591), 
        .ZN(n229) );
  OAI21_X1 U290 ( .B1(n227), .B2(n228), .A(n229), .ZN(mult_x_6_n588) );
  XNOR2_X1 U291 ( .A(mult_x_6_n1454), .B(n6901), .ZN(n230) );
  XNOR2_X1 U292 ( .A(n230), .B(mult_x_6_n727), .ZN(mult_result_w[29]) );
  INV_X1 U293 ( .A(mult_x_6_n276), .ZN(n231) );
  AOI21_X1 U294 ( .B1(n647), .B2(n648), .A(n231), .ZN(n232) );
  AOI211_X1 U295 ( .C1(n651), .C2(n655), .A(n649), .B(n232), .ZN(n233) );
  XNOR2_X1 U296 ( .A(mult_x_6_n341), .B(mult_x_6_n343), .ZN(n234) );
  XNOR2_X1 U297 ( .A(n234), .B(n233), .ZN(n235) );
  AOI22_X1 U298 ( .A1(n2580), .A2(result_o[27]), .B1(dividend_q[27]), .B2(
        n2581), .ZN(n236) );
  OAI21_X1 U299 ( .B1(n2799), .B2(n7600), .A(n236), .ZN(n237) );
  AOI21_X1 U300 ( .B1(n2571), .B2(C22_DATA3_27), .A(n237), .ZN(n238) );
  XOR2_X1 U301 ( .A(mult_x_6_n304), .B(mult_x_6_n763), .Z(n239) );
  NAND2_X1 U302 ( .A1(mult_x_6_n1456), .A2(n239), .ZN(n240) );
  OAI211_X1 U303 ( .C1(mult_x_6_n1456), .C2(n239), .A(n2579), .B(n240), .ZN(
        n241) );
  OAI211_X1 U304 ( .C1(n387), .C2(n235), .A(n238), .B(n241), .ZN(n444) );
  NAND2_X1 U305 ( .A1(result_o[17]), .A2(n2580), .ZN(n242) );
  OAI21_X1 U306 ( .B1(n8600), .B2(n2799), .A(n242), .ZN(n243) );
  AOI21_X1 U307 ( .B1(dividend_q[17]), .B2(n2581), .A(n243), .ZN(n244) );
  AOI22_X1 U308 ( .A1(C22_DATA3_17), .A2(n2571), .B1(n2579), .B2(
        mult_result_w[17]), .ZN(n245) );
  XOR2_X1 U309 ( .A(mult_x_6_n282), .B(mult_x_6_n414), .Z(n246) );
  NAND2_X1 U310 ( .A1(mult_x_6_n405), .A2(n246), .ZN(n247) );
  OAI211_X1 U311 ( .C1(mult_x_6_n405), .C2(n246), .A(n247), .B(n2578), .ZN(
        n248) );
  NAND3_X1 U312 ( .A1(n244), .A2(n245), .A3(n248), .ZN(n434) );
  INV_X1 U313 ( .A(n945), .ZN(n249) );
  NAND3_X1 U314 ( .A1(n2309), .A2(n2311), .A3(n249), .ZN(n250) );
  NOR2_X1 U315 ( .A1(n2309), .A2(n2305), .ZN(n251) );
  AOI211_X1 U316 ( .C1(n251), .C2(n945), .A(n609), .B(n2313), .ZN(n252) );
  NOR2_X1 U317 ( .A1(n609), .A2(n2578), .ZN(n253) );
  AOI21_X1 U318 ( .B1(n252), .B2(n250), .A(n253), .ZN(n447) );
  OAI21_X1 U319 ( .B1(mult_x_6_n330), .B2(mult_x_6_n1482), .A(n2579), .ZN(n254) );
  AOI21_X1 U320 ( .B1(mult_x_6_n330), .B2(mult_x_6_n1482), .A(n254), .ZN(n255)
         );
  OAI22_X1 U321 ( .A1(n2525), .A2(n2486), .B1(n2487), .B2(n2448), .ZN(n256) );
  AOI211_X1 U322 ( .C1(C22_DATA3_1), .C2(n2571), .A(n255), .B(n256), .ZN(n257)
         );
  XOR2_X1 U323 ( .A(n912), .B(mult_x_6_n647), .Z(n258) );
  NAND2_X1 U324 ( .A1(mult_x_6_n1450), .A2(n258), .ZN(n259) );
  OAI211_X1 U325 ( .C1(mult_x_6_n1450), .C2(n258), .A(n2578), .B(n259), .ZN(
        n260) );
  OAI211_X1 U326 ( .C1(n102), .C2(n2799), .A(n257), .B(n260), .ZN(n418) );
  XOR2_X1 U327 ( .A(mult_x_6_n1361), .B(mult_x_6_n787), .Z(n261) );
  XNOR2_X1 U328 ( .A(n847), .B(n261), .ZN(mult_x_6_n785) );
  INV_X1 U329 ( .A(mult_x_6_n1399), .ZN(n262) );
  INV_X1 U330 ( .A(mult_x_6_n875), .ZN(n263) );
  OAI21_X1 U331 ( .B1(mult_x_6_n875), .B2(mult_x_6_n1399), .A(mult_x_6_n884), 
        .ZN(n264) );
  OAI21_X1 U332 ( .B1(n262), .B2(n263), .A(n264), .ZN(mult_x_6_n872) );
  AOI222_X1 U333 ( .A1(mul_operand_b_q[13]), .A2(mul_operand_b_q[14]), .B1(
        mul_operand_b_q[13]), .B2(mult_x_6_n1058), .C1(mul_operand_b_q[14]), 
        .C2(mult_x_6_n1058), .ZN(n761) );
  AND2_X1 U334 ( .A1(n1010), .A2(n2196), .ZN(mult_x_6_n977) );
  INV_X1 U335 ( .A(n2173), .ZN(n265) );
  AOI21_X1 U336 ( .B1(n1010), .B2(n2196), .A(n265), .ZN(mult_x_6_n976) );
  XNOR2_X1 U337 ( .A(n2194), .B(mul_operand_b_q[4]), .ZN(n266) );
  NAND3_X1 U338 ( .A1(n2259), .A2(n2257), .A3(n2258), .ZN(n267) );
  XNOR2_X1 U339 ( .A(n267), .B(n266), .ZN(mult_x_6_n1100) );
  AOI222_X1 U340 ( .A1(mult_x_6_n693), .A2(mult_x_6_n710), .B1(mult_x_6_n693), 
        .B2(mult_x_6_n1356), .C1(mult_x_6_n710), .C2(mult_x_6_n1356), .ZN(n977) );
  INV_X1 U341 ( .A(n2364), .ZN(n268) );
  AOI21_X1 U342 ( .B1(mult_x_6_n1053), .B2(n268), .A(n2429), .ZN(n269) );
  XOR2_X1 U343 ( .A(mul_operand_b_q[19]), .B(mul_operand_b_q[20]), .Z(n270) );
  XNOR2_X1 U344 ( .A(n269), .B(n270), .ZN(mult_x_6_n1084) );
  INV_X1 U345 ( .A(n2308), .ZN(n271) );
  NOR2_X1 U346 ( .A1(n2428), .A2(n271), .ZN(n946) );
  NAND2_X1 U347 ( .A1(mult_x_6_n1078), .A2(n2225), .ZN(n272) );
  AOI222_X1 U348 ( .A1(mul_operand_b_q[25]), .A2(n608), .B1(
        mul_operand_b_q[26]), .B2(n385), .C1(n2183), .C2(n2224), .ZN(n273) );
  NAND2_X1 U349 ( .A1(n272), .A2(n273), .ZN(n274) );
  XNOR2_X1 U350 ( .A(n274), .B(n1013), .ZN(mult_x_6_n1457) );
  OAI21_X1 U351 ( .B1(n2299), .B2(n275), .A(n276), .ZN(n2303) );
  INV_X1 U352 ( .A(mult_x_6_n341), .ZN(n275) );
  INV_X1 U353 ( .A(n2302), .ZN(n276) );
  NAND2_X1 U354 ( .A1(n2225), .A2(mult_x_6_n1096), .ZN(n277) );
  AOI222_X1 U355 ( .A1(n385), .A2(mul_operand_b_q[8]), .B1(n608), .B2(
        mul_operand_b_q[7]), .C1(n2189), .C2(n2224), .ZN(n278) );
  NAND2_X1 U356 ( .A1(n278), .A2(n277), .ZN(n279) );
  XOR2_X1 U357 ( .A(mul_operand_a_q[2]), .B(n279), .Z(mult_x_6_n1475) );
  AOI222_X1 U358 ( .A1(mul_operand_b_q[8]), .A2(n608), .B1(n2186), .B2(n385), 
        .C1(mul_operand_b_q[7]), .C2(n2224), .ZN(n280) );
  NAND2_X1 U359 ( .A1(mult_x_6_n1095), .A2(n2225), .ZN(n281) );
  NAND2_X1 U360 ( .A1(n281), .A2(n280), .ZN(n282) );
  XNOR2_X1 U361 ( .A(n282), .B(n1013), .ZN(mult_x_6_n1474) );
  AOI222_X1 U362 ( .A1(n2192), .A2(n2224), .B1(n2190), .B2(n608), .C1(n2189), 
        .C2(n385), .ZN(n283) );
  NAND2_X1 U363 ( .A1(n2225), .A2(mult_x_6_n1098), .ZN(n284) );
  NAND2_X1 U364 ( .A1(n284), .A2(n283), .ZN(n285) );
  XNOR2_X1 U365 ( .A(n285), .B(n1013), .ZN(mult_x_6_n1477) );
  AOI22_X1 U366 ( .A1(n2179), .A2(n2141), .B1(n2177), .B2(n385), .ZN(n286) );
  AOI22_X1 U367 ( .A1(n2225), .A2(mult_x_6_n1072), .B1(n2224), .B2(n2180), 
        .ZN(n287) );
  NAND2_X1 U368 ( .A1(n287), .A2(n286), .ZN(n288) );
  XNOR2_X1 U369 ( .A(n288), .B(n1013), .ZN(mult_x_6_n1451) );
  AOI22_X1 U370 ( .A1(n2580), .A2(result_o[15]), .B1(dividend_q[15]), .B2(
        n2581), .ZN(n289) );
  XOR2_X1 U371 ( .A(mult_x_6_n427), .B(mult_x_6_n437), .Z(n291) );
  OAI21_X1 U372 ( .B1(n906), .B2(n291), .A(n2578), .ZN(n322) );
  AOI21_X1 U373 ( .B1(n906), .B2(n291), .A(n322), .ZN(n323) );
  XOR2_X1 U374 ( .A(mult_x_6_n1468), .B(mult_x_6_n927), .Z(n324) );
  OAI21_X1 U375 ( .B1(mult_x_6_n316), .B2(n324), .A(n2579), .ZN(n325) );
  AOI21_X1 U376 ( .B1(mult_x_6_n316), .B2(n324), .A(n325), .ZN(n326) );
  AOI211_X1 U377 ( .C1(n2571), .C2(C22_DATA3_15), .A(n323), .B(n326), .ZN(n327) );
  OAI211_X1 U378 ( .C1(n2799), .C2(n8800), .A(n289), .B(n327), .ZN(n432) );
  AOI22_X1 U379 ( .A1(n2581), .A2(dividend_q[12]), .B1(n2580), .B2(
        result_o[12]), .ZN(n328) );
  XOR2_X1 U380 ( .A(mult_x_6_n463), .B(mult_x_6_n475), .Z(n329) );
  OAI21_X1 U381 ( .B1(n2339), .B2(n643), .A(n642), .ZN(n330) );
  OAI21_X1 U382 ( .B1(n329), .B2(n330), .A(n2578), .ZN(n331) );
  AOI21_X1 U383 ( .B1(n329), .B2(n330), .A(n331), .ZN(n332) );
  XNOR2_X1 U384 ( .A(mult_x_6_n1471), .B(mult_x_6_n953), .ZN(n333) );
  OAI21_X1 U385 ( .B1(n2341), .B2(n333), .A(n2579), .ZN(n334) );
  AOI21_X1 U386 ( .B1(n2341), .B2(n333), .A(n334), .ZN(n335) );
  AOI211_X1 U387 ( .C1(n2571), .C2(C22_DATA3_12), .A(n332), .B(n335), .ZN(n336) );
  OAI211_X1 U388 ( .C1(n2799), .C2(n91), .A(n328), .B(n336), .ZN(n429) );
  OAI21_X1 U389 ( .B1(mult_x_6_n329), .B2(mult_x_6_n1481), .A(n2994), .ZN(n337) );
  AOI21_X1 U390 ( .B1(mult_x_6_n329), .B2(mult_x_6_n1481), .A(n337), .ZN(n338)
         );
  OAI22_X1 U391 ( .A1(n2447), .A2(n2487), .B1(n2527), .B2(n2486), .ZN(n339) );
  AOI211_X1 U392 ( .C1(C22_DATA3_2), .C2(n2571), .A(n338), .B(n339), .ZN(n340)
         );
  XOR2_X1 U393 ( .A(mult_x_6_n297), .B(mult_x_6_n628), .Z(n341) );
  NAND2_X1 U394 ( .A1(mult_x_6_n646), .A2(n341), .ZN(n342) );
  OAI211_X1 U395 ( .C1(mult_x_6_n646), .C2(n341), .A(n2578), .B(n342), .ZN(
        n343) );
  OAI211_X1 U396 ( .C1(n101), .C2(n2799), .A(n340), .B(n343), .ZN(n419) );
  XNOR2_X1 U397 ( .A(mult_x_6_n270), .B(n2241), .ZN(n344) );
  AOI21_X1 U398 ( .B1(C22_DATA3_29), .B2(n2571), .A(n2798), .ZN(n345) );
  NAND2_X1 U399 ( .A1(n2579), .A2(mult_result_w[29]), .ZN(n346) );
  OAI211_X1 U400 ( .C1(n387), .C2(n344), .A(n345), .B(n346), .ZN(n446) );
  XNOR2_X1 U401 ( .A(n862), .B(n866), .ZN(mult_result_w[14]) );
  XNOR2_X1 U402 ( .A(n803), .B(n804), .ZN(mult_result_w[21]) );
  XNOR2_X1 U403 ( .A(n768), .B(n769), .ZN(mult_result_w[16]) );
  XNOR2_X1 U404 ( .A(mult_x_6_n295), .B(n920), .ZN(mult_result_w[36]) );
  XNOR2_X1 U405 ( .A(n916), .B(n915), .ZN(mult_result_w[52]) );
  XNOR2_X1 U406 ( .A(mult_x_6_n292), .B(n936), .ZN(mult_result_w[39]) );
  INV_X4 U407 ( .A(n1359), .ZN(n2154) );
  BUF_X4 U408 ( .A(n2047), .Z(n2219) );
  OR2_X2 U409 ( .A1(n19601), .A2(n2049), .ZN(n2427) );
  INV_X2 U410 ( .A(n2427), .ZN(n2221) );
  INV_X4 U411 ( .A(n1774), .ZN(n2146) );
  INV_X2 U412 ( .A(n2215), .ZN(n1020) );
  INV_X4 U413 ( .A(n1149), .ZN(n2158) );
  INV_X4 U414 ( .A(n1254), .ZN(n2156) );
  INV_X4 U415 ( .A(n2574), .ZN(n2573) );
  AND2_X2 U416 ( .A1(n1671), .A2(n2147), .ZN(n1767) );
  BUF_X2 U417 ( .A(n1767), .Z(n2204) );
  INV_X4 U418 ( .A(n1569), .ZN(n2150) );
  INV_X4 U419 ( .A(n1672), .ZN(n2148) );
  NAND3_X2 U420 ( .A1(n971), .A2(n969), .A3(n966), .ZN(mult_x_6_n1098) );
  BUF_X2 U421 ( .A(mult_x_6_n1093), .Z(n2287) );
  INV_X4 U422 ( .A(mul_operand_a_q[2]), .ZN(n1013) );
  XNOR2_X1 U423 ( .A(mul_operand_b_q[8]), .B(mul_operand_b_q[7]), .ZN(n351) );
  XNOR2_X1 U424 ( .A(mult_x_6_n1439), .B(mult_x_6_n955), .ZN(n352) );
  INV_X4 U425 ( .A(n1008), .ZN(n1009) );
  INV_X1 U426 ( .A(n926), .ZN(mult_x_6_n275) );
  OAI21_X2 U427 ( .B1(n931), .B2(n2333), .A(n2409), .ZN(mult_x_6_n276) );
  BUF_X2 U428 ( .A(n1024), .Z(n355) );
  XNOR2_X1 U454 ( .A(mult_x_6_n276), .B(n925), .ZN(mult_result_w[55]) );
  OAI21_X1 U455 ( .B1(n2339), .B2(n645), .A(n644), .ZN(n641) );
  AOI21_X2 U456 ( .B1(mult_x_6_n292), .B2(n937), .A(n876), .ZN(n2339) );
  BUF_X1 U457 ( .A(n2145), .Z(n405) );
  AND2_X2 U458 ( .A1(n1148), .A2(n2157), .ZN(n1245) );
  BUF_X1 U459 ( .A(n1768), .Z(n6301) );
  AND2_X1 U460 ( .A1(n1463), .A2(n2151), .ZN(n1560) );
  INV_X2 U461 ( .A(n1464), .ZN(n2152) );
  BUF_X2 U462 ( .A(n2142), .Z(n385) );
  BUF_X1 U463 ( .A(mul_operand_b_q[5]), .Z(n2191) );
  INV_X1 U464 ( .A(n2578), .ZN(n387) );
  INV_X1 U465 ( .A(n2419), .ZN(n2202) );
  INV_X1 U466 ( .A(n2210), .ZN(n602) );
  INV_X1 U467 ( .A(n2425), .ZN(n606) );
  INV_X1 U468 ( .A(n2425), .ZN(n2203) );
  INV_X1 U469 ( .A(n2419), .ZN(n605) );
  AND3_X2 U470 ( .A1(n2159), .A2(n1059), .A3(n1060), .ZN(n2132) );
  AND2_X1 U471 ( .A1(n1358), .A2(n2153), .ZN(n1455) );
  AND2_X2 U472 ( .A1(n1568), .A2(n2149), .ZN(n1665) );
  AND2_X1 U473 ( .A1(n1253), .A2(n2155), .ZN(n1350) );
  AND2_X2 U474 ( .A1(n1060), .A2(n1142), .ZN(n2134) );
  NOR2_X1 U475 ( .A1(n1873), .A2(n1874), .ZN(n1959) );
  XNOR2_X1 U476 ( .A(n1017), .B(n1015), .ZN(mult_x_6_n1103) );
  BUF_X1 U477 ( .A(n1015), .Z(n2195) );
  AND2_X1 U478 ( .A1(n2399), .A2(mul_operand_a_q[0]), .ZN(n2142) );
  NOR2_X1 U479 ( .A1(n2428), .A2(n1000), .ZN(n999) );
  NAND2_X1 U480 ( .A1(n2428), .A2(n2308), .ZN(n998) );
  NOR2_X1 U481 ( .A1(mult_x_6_n847), .A2(mult_x_6_n1397), .ZN(n843) );
  NAND2_X2 U482 ( .A1(n2568), .A2(n2566), .ZN(n2710) );
  INV_X4 U483 ( .A(n2500), .ZN(n406) );
  AOI21_X1 U484 ( .B1(mult_x_6_n910), .B2(n722), .A(n717), .ZN(n716) );
  OR2_X1 U485 ( .A1(mult_x_6_n961), .A2(mult_x_6_n1472), .ZN(n8301) );
  NOR2_X1 U486 ( .A1(mult_x_6_n941), .A2(mult_x_6_n1405), .ZN(n2401) );
  NAND3_X1 U487 ( .A1(n2253), .A2(n2252), .A3(n2251), .ZN(mult_x_6_n1063) );
  BUF_X1 U488 ( .A(mult_x_6_n1097), .Z(n612) );
  XNOR2_X1 U489 ( .A(n696), .B(n633), .ZN(mult_x_6_n1374) );
  NOR2_X1 U490 ( .A1(n2573), .A2(n2474), .ZN(n6601) );
  BUF_X1 U491 ( .A(mult_x_6_n1100), .Z(n622) );
  INV_X1 U492 ( .A(n2418), .ZN(n627) );
  BUF_X1 U493 ( .A(n1455), .Z(n625) );
  BUF_X1 U494 ( .A(n1350), .Z(n623) );
  BUF_X1 U495 ( .A(n2144), .Z(n624) );
  INV_X1 U496 ( .A(n2417), .ZN(n626) );
  INV_X1 U497 ( .A(n2426), .ZN(n2207) );
  BUF_X1 U498 ( .A(n2145), .Z(n2226) );
  BUF_X1 U499 ( .A(n1958), .Z(n2214) );
  BUF_X1 U500 ( .A(n1561), .Z(n631) );
  BUF_X1 U501 ( .A(n1869), .Z(n629) );
  BUF_X1 U502 ( .A(n1959), .Z(n2218) );
  BUF_X1 U503 ( .A(n1868), .Z(n2209) );
  INV_X2 U504 ( .A(n2416), .ZN(n603) );
  BUF_X2 U505 ( .A(n2133), .Z(n604) );
  BUF_X2 U506 ( .A(n2119), .Z(n2224) );
  AND2_X2 U507 ( .A1(n1773), .A2(n1010), .ZN(n1868) );
  NAND2_X1 U508 ( .A1(mul_operand_b_q[27]), .A2(n2181), .ZN(n2275) );
  BUF_X2 U509 ( .A(n1456), .Z(n607) );
  BUF_X2 U510 ( .A(n2141), .Z(n608) );
  XOR2_X1 U511 ( .A(mul_operand_a_q[8]), .B(mul_operand_a_q[7]), .Z(n1874) );
  BUF_X1 U512 ( .A(mul_operand_b_q[6]), .Z(n2189) );
  XNOR2_X1 U513 ( .A(n919), .B(n918), .ZN(mult_result_w[57]) );
  INV_X1 U514 ( .A(n1003), .ZN(n1027) );
  AOI21_X1 U515 ( .B1(n641), .B2(n1004), .A(n1006), .ZN(n1003) );
  NOR2_X1 U516 ( .A1(n667), .A2(n948), .ZN(n666) );
  OAI21_X1 U517 ( .B1(n2373), .B2(n2374), .A(n2238), .ZN(n912) );
  INV_X1 U518 ( .A(n651), .ZN(n648) );
  OR2_X1 U519 ( .A1(mult_x_6_n646), .A2(mult_x_6_n628), .ZN(n944) );
  AND2_X1 U520 ( .A1(mult_x_6_n646), .A2(mult_x_6_n628), .ZN(n943) );
  INV_X1 U521 ( .A(n639), .ZN(n638) );
  NAND2_X1 U522 ( .A1(n949), .A2(n669), .ZN(n668) );
  OAI21_X1 U523 ( .B1(n654), .B2(n6501), .A(n659), .ZN(n649) );
  OAI21_X1 U524 ( .B1(n642), .B2(n942), .A(n878), .ZN(n639) );
  AOI21_X1 U525 ( .B1(n654), .B2(n653), .A(n652), .ZN(n651) );
  INV_X1 U526 ( .A(n657), .ZN(n653) );
  AND2_X1 U527 ( .A1(n2303), .A2(n950), .ZN(n949) );
  OR2_X1 U528 ( .A1(n643), .A2(n942), .ZN(n6401) );
  NAND2_X1 U529 ( .A1(n657), .A2(mult_x_6_n346), .ZN(n647) );
  INV_X1 U530 ( .A(n655), .ZN(n654) );
  OAI21_X1 U531 ( .B1(n671), .B2(n656), .A(n6701), .ZN(n655) );
  INV_X1 U532 ( .A(n671), .ZN(n669) );
  NOR2_X1 U533 ( .A1(n671), .A2(n658), .ZN(n657) );
  OR2_X1 U534 ( .A1(n645), .A2(n1002), .ZN(n643) );
  NAND2_X1 U535 ( .A1(n672), .A2(n917), .ZN(n671) );
  INV_X1 U536 ( .A(n1005), .ZN(n1002) );
  OR2_X1 U537 ( .A1(n2338), .A2(n935), .ZN(n645) );
  XNOR2_X1 U538 ( .A(mult_x_6_n706), .B(n996), .ZN(mult_x_6_n687) );
  INV_X1 U539 ( .A(n2337), .ZN(n672) );
  OAI21_X1 U540 ( .B1(n636), .B2(n635), .A(n634), .ZN(n513) );
  AND2_X1 U541 ( .A1(mult_x_6_n372), .A2(mult_x_6_n378), .ZN(n877) );
  INV_X1 U542 ( .A(n2413), .ZN(n1006) );
  OR2_X1 U543 ( .A1(mult_x_6_n340), .A2(mult_x_6_n337), .ZN(n950) );
  AND2_X1 U544 ( .A1(mult_x_6_n396), .A2(mult_x_6_n404), .ZN(n907) );
  XNOR2_X1 U545 ( .A(mult_x_6_n426), .B(mult_x_6_n415), .ZN(n898) );
  INV_X1 U546 ( .A(n2254), .ZN(n659) );
  XNOR2_X1 U547 ( .A(mult_x_6_n372), .B(mult_x_6_n378), .ZN(n930) );
  OR2_X1 U548 ( .A1(mult_x_6_n372), .A2(mult_x_6_n378), .ZN(n932) );
  AND2_X1 U549 ( .A1(mult_x_6_n571), .A2(mult_x_6_n588), .ZN(n921) );
  OR2_X1 U550 ( .A1(mult_x_6_n352), .A2(mult_x_6_n347), .ZN(n917) );
  INV_X1 U551 ( .A(n2343), .ZN(n1004) );
  NAND2_X1 U552 ( .A1(n939), .A2(n938), .ZN(n937) );
  OR2_X1 U553 ( .A1(mult_x_6_n426), .A2(mult_x_6_n415), .ZN(n902) );
  XNOR2_X1 U554 ( .A(mult_x_6_n352), .B(mult_x_6_n347), .ZN(n918) );
  OR2_X1 U555 ( .A1(mult_x_6_n571), .A2(mult_x_6_n588), .ZN(n940) );
  OR2_X1 U556 ( .A1(mult_x_6_n396), .A2(mult_x_6_n404), .ZN(n934) );
  XNOR2_X1 U557 ( .A(DP_OP_56J3_124_887_n2), .B(DP_OP_56J3_124_887_n1), .ZN(
        n636) );
  INV_X1 U558 ( .A(n927), .ZN(n658) );
  NOR2_X1 U559 ( .A1(mult_x_6_n463), .A2(mult_x_6_n475), .ZN(n942) );
  NOR2_X1 U560 ( .A1(mult_x_6_n506), .A2(mult_x_6_n520), .ZN(n935) );
  INV_X1 U561 ( .A(n886), .ZN(n656) );
  XNOR2_X1 U562 ( .A(mult_x_6_n589), .B(mult_x_6_n608), .ZN(n920) );
  INV_X1 U563 ( .A(mult_x_6_n553), .ZN(n938) );
  NAND2_X1 U564 ( .A1(mult_x_6_n727), .A2(mult_x_6_n1454), .ZN(n688) );
  XNOR2_X1 U565 ( .A(mult_x_6_n536), .B(mult_x_6_n553), .ZN(n936) );
  OR2_X1 U566 ( .A1(mult_x_6_n589), .A2(mult_x_6_n608), .ZN(n924) );
  NAND2_X1 U567 ( .A1(mult_x_6_n589), .A2(mult_x_6_n608), .ZN(n922) );
  NAND2_X1 U568 ( .A1(mult_x_6_n463), .A2(mult_x_6_n475), .ZN(n878) );
  XNOR2_X1 U569 ( .A(mult_x_6_n358), .B(mult_x_6_n363), .ZN(n925) );
  OR2_X1 U570 ( .A1(mult_x_6_n363), .A2(mult_x_6_n358), .ZN(n927) );
  XNOR2_X1 U571 ( .A(mult_x_6_n591), .B(n893), .ZN(mult_x_6_n589) );
  OR2_X1 U572 ( .A1(mult_x_6_n385), .A2(mult_x_6_n379), .ZN(n914) );
  NAND2_X1 U573 ( .A1(mult_x_6_n379), .A2(mult_x_6_n385), .ZN(n913) );
  AND2_X1 U574 ( .A1(mult_x_6_n358), .A2(mult_x_6_n363), .ZN(n886) );
  OR2_X1 U575 ( .A1(mult_x_6_n405), .A2(mult_x_6_n414), .ZN(n909) );
  INV_X1 U576 ( .A(mult_x_6_n536), .ZN(n939) );
  XNOR2_X1 U577 ( .A(mult_x_6_n379), .B(mult_x_6_n385), .ZN(n915) );
  NAND2_X1 U578 ( .A1(mult_x_6_n405), .A2(mult_x_6_n414), .ZN(n908) );
  INV_X1 U579 ( .A(mult_x_6_n346), .ZN(n6501) );
  AND2_X1 U580 ( .A1(mult_x_6_n346), .A2(mult_x_6_n344), .ZN(n2254) );
  NAND2_X1 U581 ( .A1(mult_x_6_n745), .A2(mult_x_6_n1455), .ZN(n879) );
  INV_X1 U582 ( .A(mult_x_6_n344), .ZN(n652) );
  XNOR2_X1 U583 ( .A(mult_x_6_n1415), .B(mult_x_6_n1383), .ZN(n893) );
  NAND2_X1 U584 ( .A1(mult_x_6_n781), .A2(mult_x_6_n1457), .ZN(n798) );
  XNOR2_X1 U585 ( .A(n2055), .B(n1013), .ZN(mult_x_6_n1453) );
  NOR2_X1 U586 ( .A1(mult_x_6_n729), .A2(mult_x_6_n1422), .ZN(n895) );
  NAND2_X1 U587 ( .A1(mult_x_6_n729), .A2(mult_x_6_n1422), .ZN(n894) );
  XOR2_X1 U588 ( .A(mult_x_6_n1041), .B(n2268), .Z(mult_x_6_n1073) );
  XNOR2_X1 U589 ( .A(n2064), .B(n1013), .ZN(mult_x_6_n1456) );
  NAND2_X1 U590 ( .A1(mult_x_6_n691), .A2(mult_x_6_n1388), .ZN(n882) );
  OR2_X1 U591 ( .A1(mult_x_6_n691), .A2(mult_x_6_n1388), .ZN(n884) );
  XNOR2_X1 U592 ( .A(n839), .B(n838), .ZN(mult_x_6_n1077) );
  OAI22_X1 U593 ( .A1(n977), .A2(n974), .B1(n976), .B2(n973), .ZN(
        mult_x_6_n670) );
  INV_X1 U594 ( .A(n871), .ZN(mult_x_6_n672) );
  NOR2_X1 U595 ( .A1(mult_x_6_n673), .A2(mult_x_6_n1355), .ZN(n974) );
  INV_X1 U596 ( .A(mult_x_6_n1355), .ZN(n976) );
  INV_X1 U597 ( .A(mult_x_6_n673), .ZN(n973) );
  AOI22_X1 U598 ( .A1(mult_x_6_n692), .A2(n872), .B1(mult_x_6_n675), .B2(
        mult_x_6_n1323), .ZN(n871) );
  XNOR2_X1 U599 ( .A(mult_x_6_n883), .B(mult_x_6_n1464), .ZN(n928) );
  OAI21_X1 U600 ( .B1(n849), .B2(n8501), .A(n848), .ZN(mult_x_6_n730) );
  OR2_X1 U601 ( .A1(mult_x_6_n883), .A2(mult_x_6_n1464), .ZN(n929) );
  XNOR2_X1 U602 ( .A(mult_x_6_n766), .B(n870), .ZN(mult_x_6_n749) );
  NAND2_X1 U603 ( .A1(mult_x_6_n785), .A2(mult_x_6_n1393), .ZN(n956) );
  AOI22_X1 U604 ( .A1(mult_x_6_n766), .A2(n869), .B1(mult_x_6_n1359), .B2(
        mult_x_6_n751), .ZN(n8501) );
  OR2_X1 U605 ( .A1(mult_x_6_n675), .A2(mult_x_6_n1323), .ZN(n872) );
  NAND2_X1 U606 ( .A1(mult_x_6_n733), .A2(mult_x_6_n1358), .ZN(n848) );
  NOR2_X1 U607 ( .A1(mult_x_6_n733), .A2(mult_x_6_n1358), .ZN(n849) );
  OR2_X1 U608 ( .A1(mult_x_6_n695), .A2(mult_x_6_n1324), .ZN(n841) );
  XNOR2_X1 U609 ( .A(mult_x_6_n695), .B(mult_x_6_n1324), .ZN(n842) );
  OR2_X1 U610 ( .A1(mult_x_6_n801), .A2(mult_x_6_n1394), .ZN(n797) );
  XNOR2_X1 U611 ( .A(mult_x_6_n751), .B(mult_x_6_n1359), .ZN(n870) );
  NAND2_X1 U612 ( .A1(mult_x_6_n801), .A2(mult_x_6_n1394), .ZN(n989) );
  INV_X1 U613 ( .A(n711), .ZN(mult_x_6_n674) );
  AOI22_X1 U614 ( .A1(mult_x_6_n694), .A2(n712), .B1(mult_x_6_n677), .B2(
        mult_x_6_n1291), .ZN(n711) );
  XNOR2_X1 U615 ( .A(mult_x_6_n694), .B(n713), .ZN(mult_x_6_n675) );
  OAI21_X1 U616 ( .B1(n846), .B2(n847), .A(n845), .ZN(mult_x_6_n784) );
  XNOR2_X1 U617 ( .A(mult_x_6_n750), .B(n796), .ZN(mult_x_6_n733) );
  XNOR2_X1 U618 ( .A(mult_x_6_n917), .B(mult_x_6_n1467), .ZN(n769) );
  INV_X1 U619 ( .A(n2710), .ZN(n635) );
  XNOR2_X1 U620 ( .A(mult_x_6_n884), .B(n758), .ZN(mult_x_6_n873) );
  XNOR2_X1 U621 ( .A(mult_x_6_n677), .B(mult_x_6_n1291), .ZN(n713) );
  XNOR2_X1 U622 ( .A(mult_x_6_n735), .B(mult_x_6_n1326), .ZN(n796) );
  XNOR2_X1 U623 ( .A(n773), .B(n772), .ZN(mult_x_6_n769) );
  NAND2_X1 U624 ( .A1(mult_x_6_n787), .A2(mult_x_6_n1361), .ZN(n845) );
  OAI21_X1 U625 ( .B1(n772), .B2(n771), .A(n7701), .ZN(mult_x_6_n768) );
  XNOR2_X1 U626 ( .A(mult_x_6_n714), .B(n701), .ZN(mult_x_6_n695) );
  NOR2_X1 U627 ( .A1(mult_x_6_n787), .A2(mult_x_6_n1361), .ZN(n846) );
  OR2_X1 U628 ( .A1(mult_x_6_n677), .A2(mult_x_6_n1291), .ZN(n712) );
  OR2_X1 U629 ( .A1(mult_x_6_n697), .A2(mult_x_6_n1292), .ZN(n7001) );
  XNOR2_X1 U630 ( .A(mult_x_6_n803), .B(mult_x_6_n1362), .ZN(n868) );
  XNOR2_X1 U631 ( .A(mult_x_6_n697), .B(mult_x_6_n1292), .ZN(n701) );
  XNOR2_X1 U632 ( .A(mult_x_6_n937), .B(mult_x_6_n1469), .ZN(n866) );
  XNOR2_X1 U633 ( .A(mult_x_6_n846), .B(n784), .ZN(mult_x_6_n833) );
  XNOR2_X1 U634 ( .A(mult_x_6_n802), .B(n791), .ZN(mult_x_6_n787) );
  XNOR2_X1 U635 ( .A(mult_x_6_n771), .B(n774), .ZN(n773) );
  XNOR2_X1 U636 ( .A(mult_x_6_n832), .B(n827), .ZN(mult_x_6_n817) );
  XNOR2_X1 U637 ( .A(mult_x_6_n819), .B(mult_x_6_n1363), .ZN(n827) );
  INV_X1 U638 ( .A(mult_x_6_n1328), .ZN(n774) );
  NAND2_X1 U639 ( .A1(mult_x_6_n771), .A2(mult_x_6_n1328), .ZN(n7701) );
  NOR2_X1 U640 ( .A1(mult_x_6_n771), .A2(mult_x_6_n1328), .ZN(n771) );
  XNOR2_X1 U641 ( .A(mult_x_6_n318), .B(n861), .ZN(mult_result_w[13]) );
  AOI22_X1 U642 ( .A1(n2967), .A2(dividend_q[31]), .B1(n2709), .B2(
        operand_ra_i[31]), .ZN(n634) );
  NAND2_X1 U643 ( .A1(mult_x_6_n909), .A2(mult_x_6_n1434), .ZN(n788) );
  XNOR2_X1 U644 ( .A(mult_x_6_n1054), .B(n682), .ZN(mult_x_6_n1086) );
  NOR2_X1 U645 ( .A1(mult_x_6_n909), .A2(mult_x_6_n1434), .ZN(n789) );
  XNOR2_X1 U646 ( .A(mult_x_6_n909), .B(mult_x_6_n1434), .ZN(n7901) );
  XNOR2_X1 U647 ( .A(n698), .B(n697), .ZN(mult_x_6_n803) );
  XNOR2_X1 U648 ( .A(n741), .B(n739), .ZN(mult_x_6_n819) );
  XNOR2_X1 U649 ( .A(mult_x_6_n835), .B(mult_x_6_n1364), .ZN(n784) );
  XNOR2_X1 U650 ( .A(mult_x_6_n752), .B(n681), .ZN(mult_x_6_n735) );
  XNOR2_X1 U651 ( .A(mult_x_6_n875), .B(mult_x_6_n1399), .ZN(n758) );
  XNOR2_X1 U652 ( .A(n831), .B(n832), .ZN(mult_result_w[11]) );
  OAI21_X1 U653 ( .B1(n741), .B2(n738), .A(n737), .ZN(n698) );
  XNOR2_X1 U654 ( .A(n727), .B(mult_x_6_n918), .ZN(mult_x_6_n909) );
  BUF_X2 U655 ( .A(n2741), .Z(n6101) );
  BUF_X1 U656 ( .A(n2500), .Z(n2572) );
  NAND2_X1 U657 ( .A1(mult_x_6_n919), .A2(mult_x_6_n1435), .ZN(n754) );
  NAND2_X1 U658 ( .A1(n674), .A2(n673), .ZN(mult_x_6_n918) );
  AOI22_X1 U659 ( .A1(mult_x_6_n848), .A2(n746), .B1(mult_x_6_n1332), .B2(
        mult_x_6_n837), .ZN(n741) );
  OAI21_X1 U660 ( .B1(n2314), .B2(n2315), .A(n2227), .ZN(n831) );
  XNOR2_X1 U661 ( .A(mult_x_6_n848), .B(n747), .ZN(mult_x_6_n835) );
  XNOR2_X1 U662 ( .A(mult_x_6_n737), .B(mult_x_6_n1294), .ZN(n681) );
  XNOR2_X1 U663 ( .A(mult_x_6_n789), .B(mult_x_6_n1329), .ZN(n791) );
  OR2_X1 U664 ( .A1(n2801), .A2(n2971), .ZN(n2500) );
  OAI21_X1 U665 ( .B1(n715), .B2(n716), .A(n714), .ZN(mult_x_6_n886) );
  XNOR2_X1 U666 ( .A(mult_x_6_n837), .B(mult_x_6_n1332), .ZN(n747) );
  OAI21_X1 U667 ( .B1(mult_x_6_n921), .B2(mult_x_6_n1403), .A(mult_x_6_n928), 
        .ZN(n674) );
  XNOR2_X1 U668 ( .A(n718), .B(n716), .ZN(mult_x_6_n887) );
  NAND2_X1 U669 ( .A1(mult_x_6_n929), .A2(mult_x_6_n1436), .ZN(n708) );
  XNOR2_X1 U670 ( .A(mult_x_6_n1402), .B(mult_x_6_n911), .ZN(n727) );
  XNOR2_X1 U671 ( .A(mult_x_6_n1056), .B(n822), .ZN(mult_x_6_n1088) );
  XNOR2_X1 U672 ( .A(mult_x_6_n1057), .B(n809), .ZN(mult_x_6_n1089) );
  XNOR2_X1 U673 ( .A(mult_x_6_n961), .B(mult_x_6_n1472), .ZN(n832) );
  XNOR2_X1 U674 ( .A(mult_x_6_n821), .B(n7401), .ZN(n739) );
  XNOR2_X1 U675 ( .A(mult_x_6_n910), .B(n723), .ZN(mult_x_6_n899) );
  XNOR2_X1 U676 ( .A(mult_x_6_n889), .B(n719), .ZN(n718) );
  XNOR2_X1 U677 ( .A(mult_x_6_n805), .B(mult_x_6_n1330), .ZN(n697) );
  AND2_X1 U678 ( .A1(mult_x_6_n961), .A2(mult_x_6_n1472), .ZN(n793) );
  AND2_X1 U679 ( .A1(n2567), .A2(n2615), .ZN(DP_OP_56J3_124_887_n132) );
  AND2_X2 U680 ( .A1(n2969), .A2(n2583), .ZN(n2709) );
  NOR2_X1 U681 ( .A1(mult_x_6_n889), .A2(mult_x_6_n1368), .ZN(n715) );
  NAND2_X1 U682 ( .A1(mult_x_6_n889), .A2(mult_x_6_n1368), .ZN(n714) );
  NOR2_X1 U683 ( .A1(mult_x_6_n821), .A2(mult_x_6_n1331), .ZN(n738) );
  NAND2_X1 U684 ( .A1(mult_x_6_n821), .A2(mult_x_6_n1331), .ZN(n737) );
  INV_X1 U685 ( .A(mult_x_6_n1368), .ZN(n719) );
  INV_X1 U686 ( .A(mult_x_6_n1331), .ZN(n7401) );
  BUF_X1 U687 ( .A(n2708), .Z(n2566) );
  INV_X2 U688 ( .A(n2499), .ZN(n611) );
  BUF_X1 U689 ( .A(n2708), .Z(n2567) );
  XNOR2_X1 U690 ( .A(mult_x_6_n920), .B(n745), .ZN(mult_x_6_n911) );
  NAND2_X1 U691 ( .A1(mult_x_6_n921), .A2(mult_x_6_n1403), .ZN(n673) );
  XNOR2_X1 U692 ( .A(mult_x_6_n1058), .B(n792), .ZN(mult_x_6_n1090) );
  NAND2_X1 U693 ( .A1(valid_i), .A2(n2582), .ZN(n2821) );
  AND2_X1 U694 ( .A1(mult_x_6_n901), .A2(mult_x_6_n1369), .ZN(n717) );
  XNOR2_X1 U695 ( .A(mult_x_6_n901), .B(mult_x_6_n1369), .ZN(n723) );
  NAND2_X1 U696 ( .A1(mult_x_6_n973), .A2(mult_x_6_n1474), .ZN(n748) );
  XNOR2_X1 U697 ( .A(mult_x_6_n1059), .B(n7601), .ZN(mult_x_6_n1091) );
  XNOR2_X1 U698 ( .A(mult_x_6_n954), .B(n805), .ZN(mult_x_6_n947) );
  XNOR2_X1 U699 ( .A(n892), .B(n891), .ZN(mult_x_6_n1092) );
  OAI21_X1 U700 ( .B1(n782), .B2(n781), .A(n7801), .ZN(mult_x_6_n940) );
  NAND2_X1 U701 ( .A1(mult_x_6_n1441), .A2(mult_x_6_n969), .ZN(n814) );
  NAND2_X1 U702 ( .A1(mult_x_6_n1406), .A2(mult_x_6_n949), .ZN(n806) );
  XNOR2_X1 U703 ( .A(mult_x_6_n1406), .B(mult_x_6_n949), .ZN(n805) );
  XNOR2_X1 U704 ( .A(mult_x_6_n913), .B(mult_x_6_n1370), .ZN(n745) );
  XNOR2_X1 U705 ( .A(n678), .B(mult_x_6_n325), .ZN(mult_result_w[6]) );
  NOR2_X1 U706 ( .A1(mult_x_6_n1441), .A2(mult_x_6_n969), .ZN(n815) );
  XNOR2_X1 U707 ( .A(n778), .B(n779), .ZN(mult_x_6_n963) );
  XNOR2_X1 U708 ( .A(mult_x_6_n1477), .B(mult_x_6_n987), .ZN(n678) );
  NAND2_X1 U709 ( .A1(mult_x_6_n987), .A2(mult_x_6_n1477), .ZN(n676) );
  NOR2_X1 U710 ( .A1(n662), .A2(n2707), .ZN(n661) );
  XNOR2_X1 U711 ( .A(mult_x_6_n1445), .B(n853), .ZN(mult_x_6_n987) );
  AOI21_X1 U712 ( .B1(mult_x_6_n1098), .B2(n2214), .A(n817), .ZN(n1007) );
  NAND2_X1 U713 ( .A1(mult_x_6_n1063), .A2(n2187), .ZN(n2246) );
  NOR2_X1 U714 ( .A1(mult_x_6_n1373), .A2(mult_x_6_n943), .ZN(n781) );
  NAND2_X1 U715 ( .A1(mult_x_6_n1373), .A2(mult_x_6_n943), .ZN(n7801) );
  XNOR2_X1 U716 ( .A(n854), .B(mult_x_6_n989), .ZN(n853) );
  XNOR2_X1 U717 ( .A(mult_x_6_n956), .B(n732), .ZN(mult_x_6_n949) );
  XNOR2_X1 U718 ( .A(mult_x_6_n1373), .B(mult_x_6_n943), .ZN(n783) );
  XNOR2_X1 U719 ( .A(mult_x_6_n974), .B(n874), .ZN(mult_x_6_n969) );
  XNOR2_X1 U720 ( .A(mult_x_6_n1374), .B(mult_x_6_n951), .ZN(n732) );
  XNOR2_X1 U721 ( .A(mult_x_6_n1409), .B(mult_x_6_n971), .ZN(n874) );
  XNOR2_X1 U722 ( .A(mult_x_6_n1408), .B(mult_x_6_n965), .ZN(n779) );
  NAND2_X1 U723 ( .A1(mult_x_6_n1408), .A2(mult_x_6_n965), .ZN(n775) );
  INV_X1 U724 ( .A(n663), .ZN(n662) );
  AND2_X1 U725 ( .A1(mult_x_6_n984), .A2(mult_x_6_n1411), .ZN(mult_x_6_n980)
         );
  AND2_X1 U726 ( .A1(n2393), .A2(n2395), .ZN(mult_x_6_n1064) );
  NOR2_X1 U727 ( .A1(n2583), .A2(n664), .ZN(n663) );
  AOI21_X1 U728 ( .B1(n1023), .B2(n2225), .A(n704), .ZN(n2439) );
  NAND2_X1 U729 ( .A1(mult_x_6_n1445), .A2(mult_x_6_n989), .ZN(n851) );
  NAND2_X1 U730 ( .A1(mult_x_6_n1447), .A2(mult_x_6_n994), .ZN(n965) );
  NAND2_X1 U731 ( .A1(n1861), .A2(n1862), .ZN(n696) );
  AND2_X1 U732 ( .A1(mult_x_6_n329), .A2(mult_x_6_n1481), .ZN(mult_x_6_n328)
         );
  NAND2_X1 U733 ( .A1(n2116), .A2(n705), .ZN(n704) );
  BUF_X1 U734 ( .A(mult_x_6_n1101), .Z(n833) );
  OR2_X1 U735 ( .A1(n2370), .A2(n2367), .ZN(n2371) );
  AND2_X1 U736 ( .A1(mult_x_6_n1482), .A2(mult_x_6_n330), .ZN(mult_x_6_n329)
         );
  NAND2_X1 U737 ( .A1(n2119), .A2(n2193), .ZN(n705) );
  BUF_X1 U738 ( .A(n1959), .Z(n2217) );
  BUF_X2 U739 ( .A(n2120), .Z(n2225) );
  XNOR2_X1 U740 ( .A(mul_operand_b_q[11]), .B(n349), .ZN(n891) );
  BUF_X2 U741 ( .A(n1666), .Z(n628) );
  XNOR2_X1 U742 ( .A(mul_operand_b_q[15]), .B(mul_operand_b_q[14]), .ZN(n809)
         );
  XNOR2_X1 U743 ( .A(n2182), .B(mul_operand_b_q[27]), .ZN(n838) );
  AND2_X1 U744 ( .A1(mul_operand_b_q[15]), .A2(n2185), .ZN(n8201) );
  OR2_X1 U745 ( .A1(n2185), .A2(mul_operand_b_q[15]), .ZN(n821) );
  XNOR2_X1 U746 ( .A(n2185), .B(mul_operand_b_q[15]), .ZN(n822) );
  XNOR2_X1 U747 ( .A(mul_operand_b_q[14]), .B(mul_operand_b_q[13]), .ZN(n792)
         );
  XNOR2_X1 U748 ( .A(mul_operand_b_q[18]), .B(mul_operand_b_q[17]), .ZN(n682)
         );
  BUF_X2 U749 ( .A(n2135), .Z(n632) );
  INV_X1 U750 ( .A(n2582), .ZN(n664) );
  BUF_X1 U751 ( .A(mul_operand_b_q[3]), .Z(n2194) );
  BUF_X1 U752 ( .A(mul_operand_b_q[9]), .Z(n2187) );
  NAND2_X1 U753 ( .A1(mul_operand_b_q[19]), .A2(mul_operand_b_q[20]), .ZN(
        n2414) );
  INV_X1 U754 ( .A(n2173), .ZN(n633) );
  BUF_X1 U755 ( .A(mul_operand_a_q[5]), .Z(n2175) );
  BUF_X2 U756 ( .A(mul_operand_b_q[3]), .Z(n2193) );
  INV_X1 U757 ( .A(n1017), .ZN(n1018) );
  XNOR2_X1 U758 ( .A(mul_operand_b_q[13]), .B(mul_operand_b_q[12]), .ZN(n7601)
         );
  NAND2_X1 U759 ( .A1(mul_operand_b_q[11]), .A2(mul_operand_b_q[12]), .ZN(n889) );
  NOR2_X1 U760 ( .A1(mul_operand_b_q[11]), .A2(mul_operand_b_q[12]), .ZN(n8901) );
  NAND2_X1 U761 ( .A1(n998), .A2(n2578), .ZN(n997) );
  NAND2_X2 U762 ( .A1(n2747), .A2(div_inst_q), .ZN(n2799) );
  XNOR2_X1 U763 ( .A(n2181), .B(mul_operand_b_q[29]), .ZN(n986) );
  NOR2_X1 U764 ( .A1(n2181), .A2(mul_operand_b_q[27]), .ZN(n983) );
  INV_X1 U765 ( .A(n637), .ZN(n941) );
  OAI21_X1 U766 ( .B1(n2339), .B2(n6401), .A(n638), .ZN(n637) );
  NAND2_X1 U767 ( .A1(n646), .A2(n654), .ZN(mult_x_6_n273) );
  NAND2_X1 U768 ( .A1(mult_x_6_n276), .A2(n657), .ZN(n646) );
  AOI21_X1 U769 ( .B1(mult_x_6_n276), .B2(n927), .A(n886), .ZN(n926) );
  AOI21_X1 U770 ( .B1(valid_i), .B2(n661), .A(n6601), .ZN(n1028) );
  NAND2_X1 U771 ( .A1(valid_i), .A2(n663), .ZN(n2708) );
  OAI21_X1 U772 ( .B1(n926), .B2(n2337), .A(n2412), .ZN(n919) );
  INV_X1 U773 ( .A(n665), .ZN(n947) );
  OAI21_X1 U774 ( .B1(n926), .B2(n668), .A(n666), .ZN(n665) );
  OR2_X1 U775 ( .A1(mult_x_6_n919), .A2(mult_x_6_n1435), .ZN(n756) );
  XNOR2_X1 U776 ( .A(n675), .B(mult_x_6_n928), .ZN(mult_x_6_n919) );
  XNOR2_X1 U777 ( .A(mult_x_6_n921), .B(mult_x_6_n1403), .ZN(n675) );
  NAND2_X1 U778 ( .A1(n677), .A2(n676), .ZN(mult_x_6_n324) );
  OAI21_X1 U779 ( .B1(mult_x_6_n987), .B2(mult_x_6_n1477), .A(mult_x_6_n325), 
        .ZN(n677) );
  OR2_X1 U780 ( .A1(mult_x_6_n929), .A2(mult_x_6_n1436), .ZN(n7101) );
  XNOR2_X1 U781 ( .A(n952), .B(n957), .ZN(mult_x_6_n783) );
  OAI21_X1 U782 ( .B1(n816), .B2(n815), .A(n814), .ZN(mult_x_6_n966) );
  INV_X1 U783 ( .A(n679), .ZN(mult_x_6_n734) );
  AOI22_X1 U784 ( .A1(mult_x_6_n752), .A2(n6801), .B1(mult_x_6_n737), .B2(
        mult_x_6_n1294), .ZN(n679) );
  OR2_X1 U785 ( .A1(mult_x_6_n737), .A2(mult_x_6_n1294), .ZN(n6801) );
  INV_X1 U786 ( .A(n683), .ZN(mult_x_6_n1051) );
  AOI21_X1 U787 ( .B1(mult_x_6_n1053), .B2(n2371), .A(n684), .ZN(n683) );
  INV_X1 U788 ( .A(n2372), .ZN(n684) );
  NAND2_X1 U789 ( .A1(n686), .A2(n685), .ZN(mult_x_6_n1053) );
  NAND2_X1 U790 ( .A1(mul_operand_b_q[18]), .A2(mul_operand_b_q[17]), .ZN(n685) );
  NAND2_X1 U791 ( .A1(mult_x_6_n1054), .A2(n687), .ZN(n686) );
  NAND2_X1 U792 ( .A1(n347), .A2(n350), .ZN(n687) );
  AOI22_X1 U793 ( .A1(mult_x_6_n714), .A2(n7001), .B1(mult_x_6_n697), .B2(
        mult_x_6_n1292), .ZN(n699) );
  INV_X1 U794 ( .A(n699), .ZN(mult_x_6_n694) );
  NAND2_X1 U795 ( .A1(n689), .A2(n688), .ZN(mult_x_6_n301) );
  OAI21_X1 U796 ( .B1(mult_x_6_n727), .B2(mult_x_6_n1454), .A(n6901), .ZN(n689) );
  NAND2_X1 U797 ( .A1(n8801), .A2(n879), .ZN(n6901) );
  NAND2_X1 U798 ( .A1(n692), .A2(n691), .ZN(mult_x_6_n762) );
  NAND2_X1 U799 ( .A1(mult_x_6_n765), .A2(mult_x_6_n1424), .ZN(n691) );
  OAI21_X1 U800 ( .B1(mult_x_6_n765), .B2(mult_x_6_n1424), .A(n693), .ZN(n692)
         );
  AOI22_X1 U801 ( .A1(n929), .A2(mult_x_6_n312), .B1(mult_x_6_n883), .B2(
        mult_x_6_n1464), .ZN(n2375) );
  XNOR2_X1 U802 ( .A(n694), .B(n1026), .ZN(mult_x_6_n1444) );
  NAND2_X1 U803 ( .A1(n731), .A2(n695), .ZN(n694) );
  XNOR2_X1 U804 ( .A(n759), .B(n2176), .ZN(mult_x_6_n1442) );
  NAND2_X1 U805 ( .A1(mult_x_6_n1063), .A2(mul_operand_b_q[8]), .ZN(n2245) );
  NAND2_X1 U806 ( .A1(n702), .A2(n802), .ZN(mult_x_6_n309) );
  NAND2_X1 U807 ( .A1(n703), .A2(n803), .ZN(n702) );
  OR2_X1 U808 ( .A1(mult_x_6_n857), .A2(mult_x_6_n1462), .ZN(n703) );
  XOR2_X1 U809 ( .A(mult_x_6_n1411), .B(mult_x_6_n984), .Z(mult_x_6_n981) );
  NAND2_X1 U810 ( .A1(n1863), .A2(n706), .ZN(n1864) );
  AOI21_X1 U811 ( .B1(n833), .B2(n2209), .A(n707), .ZN(n706) );
  AND2_X1 U812 ( .A1(n602), .A2(n1009), .ZN(n707) );
  INV_X1 U813 ( .A(mult_x_6_n858), .ZN(n855) );
  XNOR2_X1 U814 ( .A(mult_x_6_n849), .B(mult_x_6_n1365), .ZN(n819) );
  XNOR2_X1 U815 ( .A(mult_x_6_n860), .B(n819), .ZN(mult_x_6_n847) );
  XNOR2_X1 U816 ( .A(n757), .B(n2354), .ZN(mult_x_6_n945) );
  NOR2_X1 U817 ( .A1(mult_x_6_n953), .A2(mult_x_6_n1471), .ZN(n2340) );
  XNOR2_X1 U818 ( .A(mult_x_6_n960), .B(n352), .ZN(mult_x_6_n953) );
  NAND2_X1 U819 ( .A1(n709), .A2(n708), .ZN(mult_x_6_n926) );
  NAND2_X1 U820 ( .A1(mult_x_6_n936), .A2(n7101), .ZN(n709) );
  XNOR2_X1 U821 ( .A(mult_x_6_n712), .B(n842), .ZN(mult_x_6_n693) );
  XNOR2_X1 U822 ( .A(mult_x_6_n693), .B(mult_x_6_n1356), .ZN(n978) );
  NAND2_X1 U823 ( .A1(n1762), .A2(n7201), .ZN(n1763) );
  AOI21_X1 U824 ( .B1(n833), .B2(n2204), .A(n721), .ZN(n7201) );
  AND2_X1 U825 ( .A1(n2148), .A2(n2195), .ZN(n721) );
  AOI21_X1 U826 ( .B1(mult_x_6_n281), .B2(n934), .A(n907), .ZN(n933) );
  OAI21_X1 U827 ( .B1(n933), .B2(n2336), .A(n2411), .ZN(n916) );
  OAI21_X1 U828 ( .B1(n941), .B2(n2297), .A(n2298), .ZN(n906) );
  OAI21_X1 U829 ( .B1(n825), .B2(n824), .A(n823), .ZN(mult_x_6_n870) );
  OR2_X1 U830 ( .A1(mult_x_6_n901), .A2(mult_x_6_n1369), .ZN(n722) );
  BUF_X1 U831 ( .A(n947), .Z(n945) );
  AOI21_X1 U832 ( .B1(mult_x_6_n1098), .B2(n2219), .A(n857), .ZN(n759) );
  OAI21_X1 U833 ( .B1(n726), .B2(n725), .A(n724), .ZN(mult_x_6_n908) );
  NAND2_X1 U834 ( .A1(mult_x_6_n1402), .A2(mult_x_6_n911), .ZN(n724) );
  NOR2_X1 U835 ( .A1(mult_x_6_n1402), .A2(mult_x_6_n911), .ZN(n725) );
  INV_X1 U836 ( .A(mult_x_6_n918), .ZN(n726) );
  NAND3_X1 U837 ( .A1(n729), .A2(n2117), .A3(n728), .ZN(n2118) );
  NAND2_X1 U838 ( .A1(n2119), .A2(n1009), .ZN(n728) );
  NAND2_X1 U839 ( .A1(mult_x_6_n1100), .A2(n2225), .ZN(n729) );
  XNOR2_X1 U840 ( .A(mult_x_6_n675), .B(mult_x_6_n1323), .ZN(n873) );
  XNOR2_X1 U841 ( .A(mult_x_6_n692), .B(n873), .ZN(mult_x_6_n673) );
  XNOR2_X1 U842 ( .A(n7301), .B(n348), .ZN(mult_x_6_n1413) );
  NOR2_X1 U843 ( .A1(n1873), .A2(n1017), .ZN(n7301) );
  NAND2_X1 U844 ( .A1(n622), .A2(n2219), .ZN(n731) );
  NAND2_X1 U845 ( .A1(n734), .A2(n733), .ZN(n778) );
  NAND2_X1 U846 ( .A1(mult_x_6_n1409), .A2(mult_x_6_n971), .ZN(n733) );
  OAI21_X1 U847 ( .B1(mult_x_6_n971), .B2(mult_x_6_n1409), .A(mult_x_6_n974), 
        .ZN(n734) );
  OAI21_X1 U848 ( .B1(n735), .B2(n789), .A(n788), .ZN(mult_x_6_n906) );
  INV_X1 U849 ( .A(mult_x_6_n916), .ZN(n735) );
  NAND2_X1 U850 ( .A1(n755), .A2(n754), .ZN(mult_x_6_n916) );
  NAND2_X1 U851 ( .A1(n736), .A2(n913), .ZN(mult_x_6_n278) );
  NAND2_X1 U852 ( .A1(n916), .A2(n914), .ZN(n736) );
  OAI21_X1 U853 ( .B1(n742), .B2(n2401), .A(n867), .ZN(mult_x_6_n938) );
  INV_X1 U854 ( .A(mult_x_6_n946), .ZN(n742) );
  OAI21_X1 U855 ( .B1(n808), .B2(n807), .A(n806), .ZN(mult_x_6_n946) );
  INV_X1 U856 ( .A(n743), .ZN(mult_x_6_n910) );
  AOI22_X1 U857 ( .A1(mult_x_6_n920), .A2(n744), .B1(mult_x_6_n913), .B2(
        mult_x_6_n1370), .ZN(n743) );
  OR2_X1 U858 ( .A1(mult_x_6_n913), .A2(mult_x_6_n1370), .ZN(n744) );
  XNOR2_X1 U859 ( .A(mult_x_6_n847), .B(mult_x_6_n1397), .ZN(n844) );
  XNOR2_X1 U860 ( .A(mult_x_6_n858), .B(n844), .ZN(mult_x_6_n845) );
  OR2_X1 U861 ( .A1(mult_x_6_n837), .A2(mult_x_6_n1332), .ZN(n746) );
  XNOR2_X1 U862 ( .A(mult_x_6_n785), .B(mult_x_6_n1393), .ZN(n952) );
  NAND2_X1 U863 ( .A1(n749), .A2(n748), .ZN(mult_x_6_n321) );
  NAND2_X1 U864 ( .A1(n753), .A2(n7501), .ZN(n749) );
  NAND2_X1 U865 ( .A1(n752), .A2(n751), .ZN(n7501) );
  INV_X1 U866 ( .A(mult_x_6_n1474), .ZN(n751) );
  INV_X1 U867 ( .A(mult_x_6_n973), .ZN(n752) );
  NAND2_X1 U868 ( .A1(n2352), .A2(n2353), .ZN(n753) );
  NAND2_X1 U869 ( .A1(mult_x_6_n926), .A2(n756), .ZN(n755) );
  XNOR2_X1 U870 ( .A(mult_x_6_n861), .B(mult_x_6_n1398), .ZN(n856) );
  XNOR2_X1 U871 ( .A(n856), .B(mult_x_6_n872), .ZN(mult_x_6_n859) );
  INV_X1 U872 ( .A(n761), .ZN(mult_x_6_n1057) );
  OAI21_X1 U873 ( .B1(n764), .B2(n763), .A(n762), .ZN(mult_x_6_n1058) );
  NAND2_X1 U874 ( .A1(mul_operand_b_q[13]), .A2(mul_operand_b_q[12]), .ZN(n762) );
  NOR2_X1 U875 ( .A1(mul_operand_b_q[13]), .A2(mul_operand_b_q[12]), .ZN(n763)
         );
  INV_X1 U876 ( .A(mult_x_6_n1059), .ZN(n764) );
  OAI21_X1 U877 ( .B1(n767), .B2(n766), .A(n765), .ZN(mult_x_6_n314) );
  NAND2_X1 U878 ( .A1(mult_x_6_n917), .A2(mult_x_6_n1467), .ZN(n765) );
  NOR2_X1 U879 ( .A1(mult_x_6_n917), .A2(mult_x_6_n1467), .ZN(n766) );
  INV_X1 U880 ( .A(n768), .ZN(n767) );
  OAI21_X1 U881 ( .B1(n2361), .B2(n2362), .A(n2272), .ZN(n768) );
  XNOR2_X1 U882 ( .A(mult_x_6_n673), .B(n976), .ZN(n975) );
  XNOR2_X1 U883 ( .A(n977), .B(n975), .ZN(mult_x_6_n671) );
  INV_X1 U884 ( .A(mult_x_6_n948), .ZN(n782) );
  OAI21_X1 U885 ( .B1(n777), .B2(n776), .A(n775), .ZN(mult_x_6_n962) );
  NOR2_X1 U886 ( .A1(mult_x_6_n1408), .A2(mult_x_6_n965), .ZN(n776) );
  INV_X1 U887 ( .A(n778), .ZN(n777) );
  XNOR2_X1 U888 ( .A(mult_x_6_n948), .B(n783), .ZN(mult_x_6_n941) );
  AOI21_X1 U889 ( .B1(n831), .B2(n8301), .A(n793), .ZN(n2341) );
  OAI21_X1 U890 ( .B1(n785), .B2(n829), .A(n828), .ZN(mult_x_6_n816) );
  INV_X1 U891 ( .A(mult_x_6_n832), .ZN(n785) );
  OAI21_X1 U892 ( .B1(n818), .B2(n787), .A(n786), .ZN(mult_x_6_n832) );
  NAND2_X1 U893 ( .A1(mult_x_6_n835), .A2(mult_x_6_n1364), .ZN(n786) );
  NOR2_X1 U894 ( .A1(mult_x_6_n835), .A2(mult_x_6_n1364), .ZN(n787) );
  XNOR2_X1 U895 ( .A(mult_x_6_n916), .B(n7901), .ZN(mult_x_6_n907) );
  OAI21_X1 U896 ( .B1(n761), .B2(n812), .A(n811), .ZN(mult_x_6_n1056) );
  INV_X1 U897 ( .A(n794), .ZN(mult_x_6_n732) );
  AOI22_X1 U898 ( .A1(mult_x_6_n750), .A2(n795), .B1(mult_x_6_n735), .B2(
        mult_x_6_n1326), .ZN(n794) );
  OR2_X1 U899 ( .A1(mult_x_6_n735), .A2(mult_x_6_n1326), .ZN(n795) );
  NAND2_X1 U900 ( .A1(n2351), .A2(n2423), .ZN(n801) );
  NAND2_X1 U901 ( .A1(n990), .A2(n797), .ZN(n955) );
  NAND2_X1 U902 ( .A1(n799), .A2(n798), .ZN(mult_x_6_n304) );
  OAI21_X1 U903 ( .B1(mult_x_6_n781), .B2(mult_x_6_n1457), .A(n8001), .ZN(n799) );
  NAND2_X1 U904 ( .A1(n2348), .A2(n2260), .ZN(n8001) );
  AOI22_X1 U905 ( .A1(mult_x_6_n712), .A2(n841), .B1(mult_x_6_n695), .B2(
        mult_x_6_n1324), .ZN(n8401) );
  INV_X1 U906 ( .A(n8401), .ZN(mult_x_6_n692) );
  NAND2_X1 U907 ( .A1(mult_x_6_n857), .A2(mult_x_6_n1462), .ZN(n802) );
  OAI21_X1 U908 ( .B1(n2375), .B2(n2376), .A(n2273), .ZN(n803) );
  NOR2_X1 U909 ( .A1(mult_x_6_n1406), .A2(mult_x_6_n949), .ZN(n807) );
  INV_X1 U910 ( .A(mult_x_6_n954), .ZN(n808) );
  INV_X1 U911 ( .A(n8101), .ZN(mult_x_6_n1055) );
  AOI21_X1 U912 ( .B1(mult_x_6_n1056), .B2(n821), .A(n8201), .ZN(n8101) );
  NAND2_X1 U913 ( .A1(mul_operand_b_q[15]), .A2(mul_operand_b_q[14]), .ZN(n811) );
  NOR2_X1 U914 ( .A1(mul_operand_b_q[15]), .A2(mul_operand_b_q[14]), .ZN(n812)
         );
  INV_X1 U915 ( .A(mult_x_6_n972), .ZN(n816) );
  XNOR2_X1 U916 ( .A(n990), .B(n813), .ZN(mult_x_6_n799) );
  XNOR2_X1 U917 ( .A(mult_x_6_n801), .B(mult_x_6_n1394), .ZN(n813) );
  INV_X1 U918 ( .A(n818), .ZN(mult_x_6_n846) );
  NAND2_X1 U919 ( .A1(mult_x_6_n873), .A2(mult_x_6_n1431), .ZN(n823) );
  NOR2_X1 U920 ( .A1(mult_x_6_n873), .A2(mult_x_6_n1431), .ZN(n824) );
  INV_X1 U921 ( .A(mult_x_6_n882), .ZN(n825) );
  OAI21_X1 U922 ( .B1(n855), .B2(n843), .A(n826), .ZN(mult_x_6_n844) );
  NAND2_X1 U923 ( .A1(mult_x_6_n847), .A2(mult_x_6_n1397), .ZN(n826) );
  XNOR2_X1 U924 ( .A(n868), .B(mult_x_6_n816), .ZN(mult_x_6_n801) );
  NAND2_X1 U925 ( .A1(mult_x_6_n819), .A2(mult_x_6_n1363), .ZN(n828) );
  NOR2_X1 U926 ( .A1(mult_x_6_n819), .A2(mult_x_6_n1363), .ZN(n829) );
  NAND2_X1 U927 ( .A1(n835), .A2(n834), .ZN(mult_x_6_n1044) );
  NAND2_X1 U928 ( .A1(n2182), .A2(mul_operand_b_q[27]), .ZN(n834) );
  NAND2_X1 U929 ( .A1(n839), .A2(n836), .ZN(n835) );
  NAND2_X1 U930 ( .A1(n354), .A2(n837), .ZN(n836) );
  NAND3_X1 U931 ( .A1(n2279), .A2(n2278), .A3(n2277), .ZN(n839) );
  NAND2_X1 U932 ( .A1(n852), .A2(n851), .ZN(mult_x_6_n986) );
  OAI21_X1 U933 ( .B1(mult_x_6_n1445), .B2(mult_x_6_n989), .A(n854), .ZN(n852)
         );
  NOR2_X1 U934 ( .A1(n961), .A2(n965), .ZN(n854) );
  NAND2_X1 U935 ( .A1(n2325), .A2(n2324), .ZN(n892) );
  OAI21_X1 U936 ( .B1(n892), .B2(n8901), .A(n889), .ZN(mult_x_6_n1059) );
  NAND2_X1 U937 ( .A1(n858), .A2(n2044), .ZN(n2045) );
  AOI22_X1 U938 ( .A1(mult_x_6_n1101), .A2(n2047), .B1(n2144), .B2(n2195), 
        .ZN(n858) );
  NAND2_X1 U939 ( .A1(n8601), .A2(n859), .ZN(mult_x_6_n316) );
  NAND2_X1 U940 ( .A1(mult_x_6_n937), .A2(mult_x_6_n1469), .ZN(n859) );
  OAI21_X1 U941 ( .B1(mult_x_6_n937), .B2(mult_x_6_n1469), .A(n862), .ZN(n8601) );
  OAI21_X1 U942 ( .B1(n865), .B2(n864), .A(n863), .ZN(n862) );
  NAND2_X1 U943 ( .A1(mult_x_6_n945), .A2(mult_x_6_n1470), .ZN(n863) );
  NOR2_X1 U944 ( .A1(mult_x_6_n945), .A2(mult_x_6_n1470), .ZN(n864) );
  INV_X1 U945 ( .A(mult_x_6_n318), .ZN(n865) );
  NAND2_X1 U946 ( .A1(mult_x_6_n941), .A2(mult_x_6_n1405), .ZN(n867) );
  OR2_X1 U947 ( .A1(mult_x_6_n751), .A2(mult_x_6_n1359), .ZN(n869) );
  NAND2_X1 U948 ( .A1(n875), .A2(n2327), .ZN(mult_x_6_n842) );
  NAND2_X1 U949 ( .A1(mult_x_6_n856), .A2(n2382), .ZN(n875) );
  AND2_X1 U950 ( .A1(mult_x_6_n536), .A2(mult_x_6_n553), .ZN(n876) );
  OAI21_X1 U951 ( .B1(n2335), .B2(n2334), .A(n2410), .ZN(mult_x_6_n292) );
  XNOR2_X1 U952 ( .A(mult_x_6_n691), .B(mult_x_6_n1388), .ZN(n885) );
  XNOR2_X1 U953 ( .A(mult_x_6_n708), .B(n885), .ZN(mult_x_6_n689) );
  OAI21_X1 U954 ( .B1(mult_x_6_n745), .B2(mult_x_6_n1455), .A(n881), .ZN(n8801) );
  NAND2_X1 U955 ( .A1(n888), .A2(n887), .ZN(n881) );
  XNOR2_X1 U956 ( .A(mult_x_6_n729), .B(mult_x_6_n1422), .ZN(n897) );
  NAND2_X1 U957 ( .A1(n883), .A2(n882), .ZN(mult_x_6_n688) );
  NAND2_X1 U958 ( .A1(mult_x_6_n708), .A2(n884), .ZN(n883) );
  NAND2_X1 U959 ( .A1(mult_x_6_n763), .A2(mult_x_6_n1456), .ZN(n887) );
  OAI21_X1 U960 ( .B1(mult_x_6_n763), .B2(mult_x_6_n1456), .A(mult_x_6_n304), 
        .ZN(n888) );
  XNOR2_X1 U961 ( .A(mult_x_6_n689), .B(mult_x_6_n1420), .ZN(n996) );
  BUF_X4 U962 ( .A(mul_operand_a_q[8]), .Z(n2174) );
  INV_X1 U963 ( .A(mult_x_6_n744), .ZN(n896) );
  OAI21_X1 U964 ( .B1(n896), .B2(n895), .A(n894), .ZN(mult_x_6_n726) );
  XNOR2_X1 U965 ( .A(n897), .B(mult_x_6_n744), .ZN(mult_x_6_n727) );
  NAND2_X1 U966 ( .A1(n899), .A2(n908), .ZN(mult_x_6_n281) );
  NAND2_X1 U967 ( .A1(mult_x_6_n282), .A2(n909), .ZN(n899) );
  NAND2_X1 U968 ( .A1(n901), .A2(n900), .ZN(mult_x_6_n282) );
  NAND2_X1 U969 ( .A1(mult_x_6_n426), .A2(mult_x_6_n415), .ZN(n900) );
  NAND2_X1 U970 ( .A1(mult_x_6_n283), .A2(n902), .ZN(n901) );
  AOI21_X1 U971 ( .B1(mult_x_6_n297), .B2(n944), .A(n943), .ZN(n2332) );
  NAND2_X1 U972 ( .A1(n923), .A2(n922), .ZN(mult_x_6_n294) );
  AOI21_X1 U973 ( .B1(mult_x_6_n294), .B2(n940), .A(n921), .ZN(n2335) );
  NAND2_X1 U974 ( .A1(n904), .A2(n903), .ZN(mult_x_6_n283) );
  NAND2_X1 U975 ( .A1(mult_x_6_n427), .A2(mult_x_6_n437), .ZN(n903) );
  NAND2_X1 U976 ( .A1(n906), .A2(n905), .ZN(n904) );
  OR2_X1 U977 ( .A1(mult_x_6_n427), .A2(mult_x_6_n437), .ZN(n905) );
  NAND2_X1 U978 ( .A1(n911), .A2(n910), .ZN(mult_x_6_n297) );
  NAND2_X1 U979 ( .A1(mult_x_6_n647), .A2(mult_x_6_n1450), .ZN(n910) );
  OAI21_X1 U980 ( .B1(mult_x_6_n647), .B2(mult_x_6_n1450), .A(n912), .ZN(n911)
         );
  OAI21_X1 U981 ( .B1(n2332), .B2(n2331), .A(n2420), .ZN(mult_x_6_n295) );
  NAND2_X1 U982 ( .A1(mult_x_6_n295), .A2(n924), .ZN(n923) );
  INV_X1 U983 ( .A(n947), .ZN(mult_x_6_n270) );
  XNOR2_X2 U984 ( .A(mult_x_6_n1064), .B(n351), .ZN(mult_x_6_n1096) );
  OAI21_X1 U985 ( .B1(n988), .B2(n2422), .A(n2397), .ZN(n990) );
  NAND2_X1 U986 ( .A1(n953), .A2(n956), .ZN(mult_x_6_n782) );
  NAND2_X1 U987 ( .A1(n957), .A2(n954), .ZN(n953) );
  OR2_X1 U988 ( .A1(mult_x_6_n785), .A2(mult_x_6_n1393), .ZN(n954) );
  NAND2_X1 U989 ( .A1(n955), .A2(n989), .ZN(n957) );
  NAND3_X1 U990 ( .A1(mult_x_6_n1102), .A2(n2047), .A3(n1026), .ZN(n958) );
  NAND2_X1 U991 ( .A1(n2144), .A2(n960), .ZN(n959) );
  NOR2_X1 U992 ( .A1(n963), .A2(n1017), .ZN(n960) );
  INV_X1 U993 ( .A(n964), .ZN(n961) );
  AND2_X1 U994 ( .A1(n2046), .A2(n963), .ZN(n962) );
  INV_X1 U995 ( .A(n1026), .ZN(n963) );
  XNOR2_X1 U996 ( .A(n965), .B(n964), .ZN(mult_x_6_n991) );
  XNOR2_X1 U997 ( .A(mult_x_6_n1069), .B(n2441), .ZN(mult_x_6_n1101) );
  NAND3_X1 U998 ( .A1(n2284), .A2(n2283), .A3(n967), .ZN(n966) );
  NOR2_X1 U999 ( .A1(n1022), .A2(n968), .ZN(n967) );
  INV_X1 U1000 ( .A(n2282), .ZN(n968) );
  OR2_X1 U1001 ( .A1(n2284), .A2(n970), .ZN(n969) );
  INV_X1 U1002 ( .A(n1022), .ZN(n970) );
  NAND2_X1 U1003 ( .A1(n972), .A2(n1022), .ZN(n971) );
  NAND2_X1 U1004 ( .A1(n2283), .A2(n2282), .ZN(n972) );
  NAND2_X1 U1005 ( .A1(mult_x_6_n1067), .A2(n2192), .ZN(n2284) );
  NAND2_X1 U1006 ( .A1(mult_x_6_n1067), .A2(n2191), .ZN(n2283) );
  XNOR2_X1 U1007 ( .A(mult_x_6_n710), .B(n978), .ZN(mult_x_6_n691) );
  XNOR2_X1 U1008 ( .A(mult_x_6_n828), .B(n979), .ZN(mult_x_6_n813) );
  XNOR2_X1 U1009 ( .A(mult_x_6_n815), .B(mult_x_6_n1427), .ZN(n979) );
  XNOR2_X1 U1010 ( .A(mult_x_6_n830), .B(n2396), .ZN(mult_x_6_n815) );
  OAI21_X1 U1011 ( .B1(n982), .B2(n981), .A(n980), .ZN(mult_x_6_n812) );
  NAND2_X1 U1012 ( .A1(mult_x_6_n815), .A2(mult_x_6_n1427), .ZN(n980) );
  NOR2_X1 U1013 ( .A1(mult_x_6_n815), .A2(mult_x_6_n1427), .ZN(n981) );
  INV_X1 U1014 ( .A(mult_x_6_n828), .ZN(n982) );
  OAI21_X1 U1015 ( .B1(n984), .B2(n983), .A(n2275), .ZN(n987) );
  INV_X1 U1016 ( .A(mult_x_6_n1044), .ZN(n984) );
  XNOR2_X1 U1017 ( .A(n987), .B(n986), .ZN(mult_x_6_n1075) );
  INV_X1 U1018 ( .A(mult_x_6_n830), .ZN(n988) );
  OAI21_X1 U1019 ( .B1(n992), .B2(n991), .A(n2436), .ZN(mult_x_6_n308) );
  NOR2_X1 U1020 ( .A1(mult_x_6_n843), .A2(mult_x_6_n1461), .ZN(n991) );
  INV_X1 U1021 ( .A(mult_x_6_n309), .ZN(n992) );
  OAI21_X1 U1022 ( .B1(n995), .B2(n994), .A(n993), .ZN(mult_x_6_n686) );
  NAND2_X1 U1023 ( .A1(mult_x_6_n689), .A2(mult_x_6_n1420), .ZN(n993) );
  NOR2_X1 U1024 ( .A1(mult_x_6_n689), .A2(mult_x_6_n1420), .ZN(n994) );
  INV_X1 U1025 ( .A(mult_x_6_n706), .ZN(n995) );
  NOR2_X1 U1026 ( .A1(n2415), .A2(n1001), .ZN(n1000) );
  INV_X1 U1027 ( .A(n2308), .ZN(n1001) );
  XNOR2_X1 U1028 ( .A(n1007), .B(n2174), .ZN(mult_x_6_n1407) );
  XOR2_X1 U1029 ( .A(mul_operand_a_q[8]), .B(mul_operand_a_q[9]), .Z(n1010) );
  INV_X1 U1030 ( .A(n2375), .ZN(n1011) );
  INV_X1 U1031 ( .A(n2332), .ZN(n1012) );
  XOR2_X1 U1032 ( .A(mul_operand_a_q[2]), .B(n1014), .Z(n2399) );
  XOR2_X1 U1033 ( .A(n2121), .B(n1025), .Z(mult_x_6_n1482) );
  INV_X1 U1034 ( .A(n1021), .ZN(n1015) );
  INV_X1 U1035 ( .A(n2335), .ZN(n1016) );
  XNOR2_X1 U1036 ( .A(n2431), .B(n1013), .ZN(mult_x_6_n1483) );
  BUF_X2 U1037 ( .A(mul_operand_b_q[0]), .Z(n2196) );
  XNOR2_X1 U1038 ( .A(n1019), .B(n2174), .ZN(mult_x_6_n1410) );
  AND2_X1 U1039 ( .A1(n1956), .A2(n1957), .ZN(n1019) );
  XNOR2_X1 U1040 ( .A(n2191), .B(n2189), .ZN(n1022) );
  XOR2_X1 U1041 ( .A(mult_x_6_n1067), .B(n2285), .Z(n1023) );
  XNOR2_X1 U1042 ( .A(n1025), .B(mul_operand_a_q[3]), .ZN(n2049) );
  AND2_X1 U1043 ( .A1(mul_operand_b_q[1]), .A2(mul_operand_b_q[0]), .ZN(
        mult_x_6_n1070) );
  INV_X1 U1044 ( .A(DP_OP_56J3_124_887_n131), .ZN(n1052) );
  INV_X1 U1045 ( .A(DP_OP_56J3_124_887_n130), .ZN(n1050) );
  INV_X1 U1046 ( .A(DP_OP_56J3_124_887_n129), .ZN(n1049) );
  INV_X1 U1047 ( .A(DP_OP_56J3_124_887_n128), .ZN(n1048) );
  INV_X1 U1048 ( .A(DP_OP_56J3_124_887_n127), .ZN(n1047) );
  INV_X1 U1049 ( .A(DP_OP_56J3_124_887_n126), .ZN(n1046) );
  INV_X1 U1050 ( .A(DP_OP_56J3_124_887_n125), .ZN(n1045) );
  INV_X1 U1051 ( .A(DP_OP_56J3_124_887_n124), .ZN(n1044) );
  INV_X1 U1052 ( .A(DP_OP_56J3_124_887_n123), .ZN(n1043) );
  INV_X1 U1053 ( .A(DP_OP_56J3_124_887_n122), .ZN(n1042) );
  INV_X1 U1054 ( .A(DP_OP_56J3_124_887_n121), .ZN(n1041) );
  INV_X1 U1055 ( .A(DP_OP_56J3_124_887_n120), .ZN(n1039) );
  INV_X1 U1056 ( .A(DP_OP_56J3_124_887_n119), .ZN(n1038) );
  INV_X1 U1057 ( .A(DP_OP_56J3_124_887_n118), .ZN(n1037) );
  INV_X1 U1058 ( .A(DP_OP_56J3_124_887_n117), .ZN(n1036) );
  INV_X1 U1059 ( .A(DP_OP_56J3_124_887_n116), .ZN(n1035) );
  INV_X1 U1060 ( .A(DP_OP_56J3_124_887_n115), .ZN(n1034) );
  INV_X1 U1061 ( .A(DP_OP_56J3_124_887_n114), .ZN(n1033) );
  INV_X1 U1062 ( .A(DP_OP_56J3_124_887_n113), .ZN(n1032) );
  INV_X1 U1063 ( .A(DP_OP_56J3_124_887_n112), .ZN(n1031) );
  INV_X1 U1064 ( .A(DP_OP_56J3_124_887_n111), .ZN(n1030) );
  INV_X1 U1065 ( .A(DP_OP_56J3_124_887_n110), .ZN(n1058) );
  INV_X1 U1066 ( .A(DP_OP_56J3_124_887_n109), .ZN(n1057) );
  INV_X1 U1067 ( .A(DP_OP_56J3_124_887_n108), .ZN(n1056) );
  INV_X1 U1068 ( .A(DP_OP_56J3_124_887_n107), .ZN(n1055) );
  INV_X1 U1069 ( .A(DP_OP_56J3_124_887_n106), .ZN(n1054) );
  INV_X1 U1070 ( .A(DP_OP_56J3_124_887_n105), .ZN(n1053) );
  INV_X1 U1071 ( .A(DP_OP_56J3_124_887_n104), .ZN(n1051) );
  INV_X1 U1072 ( .A(DP_OP_56J3_124_887_n103), .ZN(n1040) );
  INV_X1 U1073 ( .A(DP_OP_56J3_124_887_n102), .ZN(n1029) );
  XOR2_X1 U1074 ( .A(mul_operand_a_q[32]), .B(mul_operand_a_q[31]), .Z(n1060)
         );
  XOR2_X1 U1075 ( .A(mul_operand_a_q[30]), .B(mul_operand_a_q[29]), .Z(n1142)
         );
  NOR2_X1 U1076 ( .A1(n1060), .A2(n2159), .ZN(n2133) );
  XNOR2_X1 U1077 ( .A(mul_operand_a_q[31]), .B(mul_operand_a_q[30]), .ZN(n1059) );
  NOR2_X1 U1078 ( .A1(n1142), .A2(n1059), .ZN(n2135) );
  AOI22_X1 U1079 ( .A1(mul_operand_b_q[32]), .A2(n604), .B1(n632), .B2(n2179), 
        .ZN(n1062) );
  AOI22_X1 U1080 ( .A1(n2132), .A2(n2180), .B1(n2134), .B2(mult_x_6_n1072), 
        .ZN(n1061) );
  NAND2_X1 U1081 ( .A1(n1062), .A2(n1061), .ZN(n2122) );
  AOI22_X1 U1082 ( .A1(n604), .A2(n2179), .B1(n632), .B2(n2180), .ZN(n1064) );
  AOI22_X1 U1083 ( .A1(n2132), .A2(mul_operand_b_q[29]), .B1(n2134), .B2(
        mult_x_6_n1073), .ZN(n1063) );
  NAND2_X1 U1084 ( .A1(n1064), .A2(n1063), .ZN(n1065) );
  XOR2_X1 U1085 ( .A(mul_operand_a_q[32]), .B(n1065), .Z(mult_x_6_n1106) );
  AOI22_X1 U1086 ( .A1(n604), .A2(n2180), .B1(n632), .B2(mul_operand_b_q[29]), 
        .ZN(n1067) );
  AOI22_X1 U1087 ( .A1(n2132), .A2(mul_operand_b_q[28]), .B1(n2134), .B2(
        mult_x_6_n1074), .ZN(n1066) );
  NAND2_X1 U1088 ( .A1(n1067), .A2(n1066), .ZN(n1068) );
  XOR2_X1 U1089 ( .A(mul_operand_a_q[32]), .B(n1068), .Z(mult_x_6_n1107) );
  AOI22_X1 U1090 ( .A1(n604), .A2(mul_operand_b_q[29]), .B1(n632), .B2(
        mul_operand_b_q[28]), .ZN(n1070) );
  AOI22_X1 U1091 ( .A1(n2132), .A2(mul_operand_b_q[27]), .B1(n2134), .B2(
        mult_x_6_n1075), .ZN(n1069) );
  NAND2_X1 U1092 ( .A1(n1070), .A2(n1069), .ZN(n1071) );
  XOR2_X1 U1093 ( .A(mul_operand_a_q[32]), .B(n1071), .Z(mult_x_6_n1108) );
  AOI22_X1 U1094 ( .A1(n604), .A2(mul_operand_b_q[28]), .B1(n632), .B2(
        mul_operand_b_q[27]), .ZN(n1073) );
  AOI22_X1 U1095 ( .A1(n2132), .A2(mul_operand_b_q[26]), .B1(n2134), .B2(
        mult_x_6_n1076), .ZN(n1072) );
  NAND2_X1 U1096 ( .A1(n1073), .A2(n1072), .ZN(n1074) );
  XOR2_X1 U1097 ( .A(mul_operand_a_q[32]), .B(n1074), .Z(mult_x_6_n1109) );
  AOI22_X1 U1098 ( .A1(n604), .A2(mul_operand_b_q[27]), .B1(n632), .B2(
        mul_operand_b_q[26]), .ZN(n1076) );
  AOI22_X1 U1099 ( .A1(n2132), .A2(mul_operand_b_q[25]), .B1(n2134), .B2(
        mult_x_6_n1077), .ZN(n1075) );
  NAND2_X1 U1100 ( .A1(n1076), .A2(n1075), .ZN(n1077) );
  XOR2_X1 U1101 ( .A(mul_operand_a_q[32]), .B(n1077), .Z(mult_x_6_n1110) );
  AOI22_X1 U1102 ( .A1(n604), .A2(mul_operand_b_q[25]), .B1(n632), .B2(
        mul_operand_b_q[24]), .ZN(n1079) );
  AOI22_X1 U1103 ( .A1(n2132), .A2(mul_operand_b_q[23]), .B1(n2134), .B2(
        mult_x_6_n1079), .ZN(n1078) );
  NAND2_X1 U1104 ( .A1(n1079), .A2(n1078), .ZN(n1080) );
  XOR2_X1 U1105 ( .A(mul_operand_a_q[32]), .B(n1080), .Z(mult_x_6_n1111) );
  AOI22_X1 U1106 ( .A1(n604), .A2(mul_operand_b_q[24]), .B1(n632), .B2(
        mul_operand_b_q[23]), .ZN(n1082) );
  AOI22_X1 U1107 ( .A1(n2132), .A2(mul_operand_b_q[22]), .B1(n2134), .B2(
        mult_x_6_n1080), .ZN(n1081) );
  NAND2_X1 U1108 ( .A1(n1082), .A2(n1081), .ZN(n1083) );
  XOR2_X1 U1109 ( .A(mul_operand_a_q[32]), .B(n1083), .Z(mult_x_6_n1112) );
  AOI22_X1 U1110 ( .A1(n604), .A2(mul_operand_b_q[23]), .B1(n632), .B2(
        mul_operand_b_q[22]), .ZN(n1085) );
  AOI22_X1 U1111 ( .A1(n2132), .A2(mul_operand_b_q[21]), .B1(n2134), .B2(
        mult_x_6_n1081), .ZN(n1084) );
  NAND2_X1 U1112 ( .A1(n1085), .A2(n1084), .ZN(n1086) );
  XOR2_X1 U1113 ( .A(mul_operand_a_q[32]), .B(n1086), .Z(mult_x_6_n1113) );
  AOI22_X1 U1114 ( .A1(n604), .A2(mul_operand_b_q[22]), .B1(n2132), .B2(
        mul_operand_b_q[20]), .ZN(n1088) );
  AOI22_X1 U1115 ( .A1(n632), .A2(mul_operand_b_q[21]), .B1(n2134), .B2(
        mult_x_6_n1082), .ZN(n1087) );
  NAND2_X1 U1116 ( .A1(n1088), .A2(n1087), .ZN(n1089) );
  XOR2_X1 U1117 ( .A(mul_operand_a_q[32]), .B(n1089), .Z(mult_x_6_n1114) );
  AOI22_X1 U1118 ( .A1(n604), .A2(mul_operand_b_q[21]), .B1(n2132), .B2(
        mul_operand_b_q[19]), .ZN(n1091) );
  AOI22_X1 U1119 ( .A1(n632), .A2(mul_operand_b_q[20]), .B1(n2134), .B2(
        mult_x_6_n1083), .ZN(n1090) );
  NAND2_X1 U1120 ( .A1(n1091), .A2(n1090), .ZN(n1092) );
  XOR2_X1 U1121 ( .A(mul_operand_a_q[32]), .B(n1092), .Z(mult_x_6_n1115) );
  AOI22_X1 U1122 ( .A1(n604), .A2(mul_operand_b_q[19]), .B1(n2132), .B2(
        mul_operand_b_q[17]), .ZN(n1094) );
  AOI22_X1 U1123 ( .A1(n632), .A2(mul_operand_b_q[18]), .B1(n2134), .B2(
        mult_x_6_n1085), .ZN(n1093) );
  NAND2_X1 U1124 ( .A1(n1094), .A2(n1093), .ZN(n1095) );
  XOR2_X1 U1125 ( .A(mul_operand_a_q[32]), .B(n1095), .Z(mult_x_6_n1116) );
  AOI22_X1 U1126 ( .A1(n604), .A2(mul_operand_b_q[18]), .B1(n2132), .B2(n2184), 
        .ZN(n1097) );
  AOI22_X1 U1127 ( .A1(n632), .A2(mul_operand_b_q[17]), .B1(n2134), .B2(
        mult_x_6_n1086), .ZN(n1096) );
  NAND2_X1 U1128 ( .A1(n1097), .A2(n1096), .ZN(n1098) );
  XOR2_X1 U1129 ( .A(mul_operand_a_q[32]), .B(n1098), .Z(mult_x_6_n1117) );
  AOI22_X1 U1130 ( .A1(n604), .A2(mul_operand_b_q[17]), .B1(n2132), .B2(
        mul_operand_b_q[15]), .ZN(n1100) );
  AOI22_X1 U1131 ( .A1(n632), .A2(n2184), .B1(n2134), .B2(mult_x_6_n1087), 
        .ZN(n1099) );
  NAND2_X1 U1132 ( .A1(n1100), .A2(n1099), .ZN(n1101) );
  XOR2_X1 U1133 ( .A(mul_operand_a_q[32]), .B(n1101), .Z(mult_x_6_n1118) );
  AOI22_X1 U1134 ( .A1(n604), .A2(n2184), .B1(n2132), .B2(mul_operand_b_q[14]), 
        .ZN(n1103) );
  AOI22_X1 U1135 ( .A1(n632), .A2(mul_operand_b_q[15]), .B1(n2134), .B2(
        mult_x_6_n1088), .ZN(n1102) );
  NAND2_X1 U1136 ( .A1(n1103), .A2(n1102), .ZN(n1104) );
  XOR2_X1 U1137 ( .A(mul_operand_a_q[32]), .B(n1104), .Z(mult_x_6_n1119) );
  AOI22_X1 U1138 ( .A1(n604), .A2(mul_operand_b_q[15]), .B1(n2132), .B2(
        mul_operand_b_q[13]), .ZN(n1106) );
  AOI22_X1 U1139 ( .A1(n632), .A2(mul_operand_b_q[14]), .B1(n2134), .B2(
        mult_x_6_n1089), .ZN(n1105) );
  NAND2_X1 U1140 ( .A1(n1106), .A2(n1105), .ZN(n1107) );
  XOR2_X1 U1141 ( .A(mul_operand_a_q[32]), .B(n1107), .Z(mult_x_6_n1120) );
  AOI22_X1 U1142 ( .A1(n604), .A2(mul_operand_b_q[13]), .B1(n2132), .B2(
        mul_operand_b_q[11]), .ZN(n1109) );
  AOI22_X1 U1143 ( .A1(n632), .A2(mul_operand_b_q[12]), .B1(n2134), .B2(
        mult_x_6_n1091), .ZN(n1108) );
  NAND2_X1 U1144 ( .A1(n1109), .A2(n1108), .ZN(n1110) );
  XOR2_X1 U1145 ( .A(mul_operand_a_q[32]), .B(n1110), .Z(mult_x_6_n1121) );
  AOI22_X1 U1146 ( .A1(n604), .A2(mul_operand_b_q[12]), .B1(n632), .B2(
        mul_operand_b_q[11]), .ZN(n1112) );
  AOI22_X1 U1147 ( .A1(n2132), .A2(mul_operand_b_q[10]), .B1(n2134), .B2(
        mult_x_6_n1092), .ZN(n1111) );
  NAND2_X1 U1148 ( .A1(n1112), .A2(n1111), .ZN(n1113) );
  XOR2_X1 U1149 ( .A(mul_operand_a_q[32]), .B(n1113), .Z(mult_x_6_n1122) );
  AOI22_X1 U1150 ( .A1(n604), .A2(mul_operand_b_q[11]), .B1(n632), .B2(
        mul_operand_b_q[10]), .ZN(n1115) );
  AOI22_X1 U1151 ( .A1(n2132), .A2(n2186), .B1(n2134), .B2(n2287), .ZN(n1114)
         );
  NAND2_X1 U1152 ( .A1(n1115), .A2(n1114), .ZN(n1116) );
  XOR2_X1 U1153 ( .A(mul_operand_a_q[32]), .B(n1116), .Z(mult_x_6_n1123) );
  AOI22_X1 U1154 ( .A1(n604), .A2(mul_operand_b_q[10]), .B1(n2132), .B2(
        mul_operand_b_q[8]), .ZN(n1118) );
  AOI22_X1 U1155 ( .A1(n632), .A2(n2186), .B1(n2134), .B2(mult_x_6_n1094), 
        .ZN(n1117) );
  NAND2_X1 U1156 ( .A1(n1118), .A2(n1117), .ZN(n1119) );
  XOR2_X1 U1157 ( .A(mul_operand_a_q[32]), .B(n1119), .Z(mult_x_6_n1124) );
  AOI22_X1 U1158 ( .A1(n604), .A2(n2186), .B1(n2132), .B2(mul_operand_b_q[7]), 
        .ZN(n1121) );
  AOI22_X1 U1159 ( .A1(n632), .A2(mul_operand_b_q[8]), .B1(n2134), .B2(
        mult_x_6_n1095), .ZN(n1120) );
  NAND2_X1 U1160 ( .A1(n1121), .A2(n1120), .ZN(n1122) );
  XOR2_X1 U1161 ( .A(mul_operand_a_q[32]), .B(n1122), .Z(mult_x_6_n1125) );
  AOI22_X1 U1162 ( .A1(n604), .A2(mul_operand_b_q[7]), .B1(n2132), .B2(n2190), 
        .ZN(n1124) );
  AOI22_X1 U1163 ( .A1(n632), .A2(n2189), .B1(n2134), .B2(n612), .ZN(n1123) );
  NAND2_X1 U1164 ( .A1(n1124), .A2(n1123), .ZN(n1125) );
  XOR2_X1 U1165 ( .A(mul_operand_a_q[32]), .B(n1125), .Z(mult_x_6_n1126) );
  AOI22_X1 U1166 ( .A1(n604), .A2(n2189), .B1(n2132), .B2(n2192), .ZN(n1127)
         );
  AOI22_X1 U1167 ( .A1(n632), .A2(n2190), .B1(n2134), .B2(mult_x_6_n1098), 
        .ZN(n1126) );
  NAND2_X1 U1168 ( .A1(n1127), .A2(n1126), .ZN(n1128) );
  XOR2_X1 U1169 ( .A(mul_operand_a_q[32]), .B(n1128), .Z(mult_x_6_n1127) );
  AOI22_X1 U1170 ( .A1(n604), .A2(n2190), .B1(n2132), .B2(n2193), .ZN(n1130)
         );
  AOI22_X1 U1171 ( .A1(n632), .A2(n2192), .B1(n2134), .B2(n355), .ZN(n1129) );
  NAND2_X1 U1172 ( .A1(n1130), .A2(n1129), .ZN(n1131) );
  XOR2_X1 U1173 ( .A(mul_operand_a_q[32]), .B(n1131), .Z(mult_x_6_n1128) );
  AOI22_X1 U1174 ( .A1(n604), .A2(n2192), .B1(n2132), .B2(n1009), .ZN(n1133)
         );
  AOI22_X1 U1175 ( .A1(n632), .A2(n2193), .B1(n2134), .B2(n622), .ZN(n1132) );
  NAND2_X1 U1176 ( .A1(n1133), .A2(n1132), .ZN(n1134) );
  XOR2_X1 U1177 ( .A(mul_operand_a_q[32]), .B(n1134), .Z(mult_x_6_n1129) );
  AOI22_X1 U1178 ( .A1(n604), .A2(n2193), .B1(n2132), .B2(n2195), .ZN(n1136)
         );
  AOI22_X1 U1179 ( .A1(n632), .A2(n1009), .B1(n833), .B2(n2134), .ZN(n1135) );
  NAND2_X1 U1180 ( .A1(n1136), .A2(n1135), .ZN(n1137) );
  XOR2_X1 U1181 ( .A(mul_operand_a_q[32]), .B(n1137), .Z(mult_x_6_n1130) );
  AOI22_X1 U1182 ( .A1(n604), .A2(n1009), .B1(n2132), .B2(n1018), .ZN(n1139)
         );
  AOI22_X1 U1183 ( .A1(n632), .A2(n2195), .B1(mult_x_6_n1102), .B2(n2134), 
        .ZN(n1138) );
  NAND2_X1 U1184 ( .A1(n1139), .A2(n1138), .ZN(n1140) );
  XOR2_X1 U1185 ( .A(mul_operand_a_q[32]), .B(n1140), .Z(mult_x_6_n1131) );
  AOI222_X1 U1186 ( .A1(n2133), .A2(n2195), .B1(n2135), .B2(n1018), .C1(n2134), 
        .C2(mult_x_6_n1103), .ZN(n1141) );
  XNOR2_X1 U1187 ( .A(mul_operand_a_q[32]), .B(n1141), .ZN(mult_x_6_n1132) );
  NAND2_X1 U1188 ( .A1(n1018), .A2(n1142), .ZN(n1143) );
  XNOR2_X1 U1189 ( .A(n1143), .B(mul_operand_a_q[32]), .ZN(mult_x_6_n1133) );
  XNOR2_X1 U1190 ( .A(mul_operand_a_q[26]), .B(mul_operand_a_q[27]), .ZN(n1147) );
  XOR2_X1 U1191 ( .A(mul_operand_a_q[29]), .B(mul_operand_a_q[28]), .Z(n1148)
         );
  XNOR2_X1 U1192 ( .A(mul_operand_a_q[28]), .B(mul_operand_a_q[27]), .ZN(n1144) );
  NAND3_X1 U1193 ( .A1(n1148), .A2(n1147), .A3(n1144), .ZN(n1149) );
  NAND3_X1 U1194 ( .A1(n1147), .A2(n1149), .A3(n2416), .ZN(n1145) );
  NAND2_X1 U1195 ( .A1(n1145), .A2(n2177), .ZN(n1146) );
  XOR2_X1 U1196 ( .A(mul_operand_a_q[29]), .B(n1146), .Z(mult_x_6_n1134) );
  NOR2_X1 U1197 ( .A1(n1147), .A2(n1148), .ZN(n1246) );
  OR2_X1 U1198 ( .A1(n1246), .A2(n603), .ZN(n1150) );
  AOI222_X1 U1199 ( .A1(n1150), .A2(mul_operand_b_q[32]), .B1(mult_x_6_n1071), 
        .B2(n1245), .C1(mul_operand_b_q[31]), .C2(n2158), .ZN(n1151) );
  XNOR2_X1 U1200 ( .A(mul_operand_a_q[29]), .B(n1151), .ZN(mult_x_6_n1135) );
  AOI22_X1 U1201 ( .A1(n2180), .A2(n2158), .B1(mult_x_6_n1072), .B2(n1245), 
        .ZN(n1153) );
  NAND2_X1 U1202 ( .A1(n2177), .A2(n1246), .ZN(n1152) );
  OAI211_X1 U1203 ( .C1(n2178), .C2(n2416), .A(n1153), .B(n1152), .ZN(n1154)
         );
  XOR2_X1 U1204 ( .A(mul_operand_a_q[29]), .B(n1154), .Z(mult_x_6_n1136) );
  AOI22_X1 U1205 ( .A1(n2179), .A2(n1246), .B1(n2180), .B2(n603), .ZN(n1156)
         );
  AOI22_X1 U1206 ( .A1(mul_operand_b_q[29]), .A2(n2158), .B1(mult_x_6_n1073), 
        .B2(n1245), .ZN(n1155) );
  NAND2_X1 U1207 ( .A1(n1156), .A2(n1155), .ZN(n1157) );
  XOR2_X1 U1208 ( .A(mul_operand_a_q[29]), .B(n1157), .Z(mult_x_6_n1137) );
  AOI22_X1 U1209 ( .A1(n2180), .A2(n1246), .B1(mul_operand_b_q[29]), .B2(n603), 
        .ZN(n1159) );
  AOI22_X1 U1210 ( .A1(n2181), .A2(n2158), .B1(mult_x_6_n1074), .B2(n1245), 
        .ZN(n1158) );
  NAND2_X1 U1211 ( .A1(n1159), .A2(n1158), .ZN(n1160) );
  XOR2_X1 U1212 ( .A(mul_operand_a_q[29]), .B(n1160), .Z(mult_x_6_n1138) );
  AOI22_X1 U1213 ( .A1(mul_operand_b_q[29]), .A2(n1246), .B1(
        mul_operand_b_q[28]), .B2(n603), .ZN(n1162) );
  AOI22_X1 U1214 ( .A1(mul_operand_b_q[27]), .A2(n2158), .B1(mult_x_6_n1075), 
        .B2(n1245), .ZN(n1161) );
  NAND2_X1 U1215 ( .A1(n1162), .A2(n1161), .ZN(n1163) );
  XOR2_X1 U1216 ( .A(mul_operand_a_q[29]), .B(n1163), .Z(mult_x_6_n1139) );
  AOI22_X1 U1217 ( .A1(n2181), .A2(n2197), .B1(mul_operand_b_q[27]), .B2(n603), 
        .ZN(n1165) );
  AOI22_X1 U1218 ( .A1(n2182), .A2(n2158), .B1(mult_x_6_n1076), .B2(n1245), 
        .ZN(n1164) );
  NAND2_X1 U1219 ( .A1(n1165), .A2(n1164), .ZN(n1166) );
  XOR2_X1 U1220 ( .A(mul_operand_a_q[29]), .B(n1166), .Z(mult_x_6_n1140) );
  AOI22_X1 U1221 ( .A1(mul_operand_b_q[27]), .A2(n2197), .B1(
        mul_operand_b_q[26]), .B2(n603), .ZN(n1168) );
  AOI22_X1 U1222 ( .A1(mul_operand_b_q[25]), .A2(n2158), .B1(mult_x_6_n1077), 
        .B2(n1245), .ZN(n1167) );
  NAND2_X1 U1223 ( .A1(n1168), .A2(n1167), .ZN(n1169) );
  XOR2_X1 U1224 ( .A(mul_operand_a_q[29]), .B(n1169), .Z(mult_x_6_n1141) );
  AOI22_X1 U1225 ( .A1(n2182), .A2(n2197), .B1(mul_operand_b_q[25]), .B2(n603), 
        .ZN(n1171) );
  AOI22_X1 U1226 ( .A1(n2183), .A2(n2158), .B1(n1245), .B2(mult_x_6_n1078), 
        .ZN(n1170) );
  NAND2_X1 U1227 ( .A1(n1171), .A2(n1170), .ZN(n1172) );
  XOR2_X1 U1228 ( .A(mul_operand_a_q[29]), .B(n1172), .Z(mult_x_6_n1142) );
  AOI22_X1 U1229 ( .A1(mul_operand_b_q[25]), .A2(n2197), .B1(
        mul_operand_b_q[24]), .B2(n603), .ZN(n1174) );
  AOI22_X1 U1230 ( .A1(mul_operand_b_q[23]), .A2(n2158), .B1(mult_x_6_n1079), 
        .B2(n1245), .ZN(n1173) );
  NAND2_X1 U1231 ( .A1(n1174), .A2(n1173), .ZN(n1175) );
  XOR2_X1 U1232 ( .A(mul_operand_a_q[29]), .B(n1175), .Z(mult_x_6_n1143) );
  AOI22_X1 U1233 ( .A1(n2183), .A2(n2197), .B1(mul_operand_b_q[23]), .B2(n603), 
        .ZN(n1177) );
  AOI22_X1 U1234 ( .A1(mul_operand_b_q[22]), .A2(n2158), .B1(mult_x_6_n1080), 
        .B2(n1245), .ZN(n1176) );
  NAND2_X1 U1235 ( .A1(n1177), .A2(n1176), .ZN(n1178) );
  XOR2_X1 U1236 ( .A(mul_operand_a_q[29]), .B(n1178), .Z(mult_x_6_n1144) );
  AOI22_X1 U1237 ( .A1(mul_operand_b_q[23]), .A2(n2197), .B1(
        mul_operand_b_q[22]), .B2(n603), .ZN(n1180) );
  AOI22_X1 U1238 ( .A1(mul_operand_b_q[21]), .A2(n2158), .B1(mult_x_6_n1081), 
        .B2(n1245), .ZN(n1179) );
  NAND2_X1 U1239 ( .A1(n1180), .A2(n1179), .ZN(n1181) );
  XOR2_X1 U1240 ( .A(mul_operand_a_q[29]), .B(n1181), .Z(mult_x_6_n1145) );
  AOI22_X1 U1241 ( .A1(mul_operand_b_q[22]), .A2(n2197), .B1(
        mul_operand_b_q[21]), .B2(n603), .ZN(n1183) );
  AOI22_X1 U1242 ( .A1(mul_operand_b_q[20]), .A2(n2158), .B1(mult_x_6_n1082), 
        .B2(n1245), .ZN(n1182) );
  NAND2_X1 U1243 ( .A1(n1183), .A2(n1182), .ZN(n1184) );
  XOR2_X1 U1244 ( .A(mul_operand_a_q[29]), .B(n1184), .Z(mult_x_6_n1146) );
  AOI22_X1 U1245 ( .A1(mul_operand_b_q[21]), .A2(n2197), .B1(
        mul_operand_b_q[20]), .B2(n603), .ZN(n1186) );
  AOI22_X1 U1246 ( .A1(mul_operand_b_q[19]), .A2(n2158), .B1(mult_x_6_n1083), 
        .B2(n1245), .ZN(n1185) );
  NAND2_X1 U1247 ( .A1(n1186), .A2(n1185), .ZN(n1187) );
  XOR2_X1 U1248 ( .A(mul_operand_a_q[29]), .B(n1187), .Z(mult_x_6_n1147) );
  AOI22_X1 U1249 ( .A1(mul_operand_b_q[20]), .A2(n2197), .B1(
        mul_operand_b_q[19]), .B2(n603), .ZN(n1189) );
  AOI22_X1 U1250 ( .A1(mul_operand_b_q[18]), .A2(n2158), .B1(n1245), .B2(
        mult_x_6_n1084), .ZN(n1188) );
  NAND2_X1 U1251 ( .A1(n1189), .A2(n1188), .ZN(n1190) );
  XOR2_X1 U1252 ( .A(mul_operand_a_q[29]), .B(n1190), .Z(mult_x_6_n1148) );
  AOI22_X1 U1253 ( .A1(mul_operand_b_q[19]), .A2(n2197), .B1(
        mul_operand_b_q[18]), .B2(n603), .ZN(n1192) );
  AOI22_X1 U1254 ( .A1(mul_operand_b_q[17]), .A2(n2158), .B1(mult_x_6_n1085), 
        .B2(n1245), .ZN(n1191) );
  NAND2_X1 U1255 ( .A1(n1192), .A2(n1191), .ZN(n1193) );
  XOR2_X1 U1256 ( .A(mul_operand_a_q[29]), .B(n1193), .Z(mult_x_6_n1149) );
  AOI22_X1 U1257 ( .A1(mul_operand_b_q[17]), .A2(n603), .B1(
        mul_operand_b_q[18]), .B2(n1246), .ZN(n1195) );
  AOI22_X1 U1258 ( .A1(n2185), .A2(n2158), .B1(mult_x_6_n1086), .B2(n1245), 
        .ZN(n1194) );
  NAND2_X1 U1259 ( .A1(n1195), .A2(n1194), .ZN(n1196) );
  XOR2_X1 U1260 ( .A(mul_operand_a_q[29]), .B(n1196), .Z(mult_x_6_n1150) );
  AOI22_X1 U1261 ( .A1(mul_operand_b_q[17]), .A2(n2197), .B1(n2184), .B2(n603), 
        .ZN(n1198) );
  AOI22_X1 U1262 ( .A1(mul_operand_b_q[15]), .A2(n2158), .B1(mult_x_6_n1087), 
        .B2(n1245), .ZN(n1197) );
  NAND2_X1 U1263 ( .A1(n1198), .A2(n1197), .ZN(n1199) );
  XOR2_X1 U1264 ( .A(mul_operand_a_q[29]), .B(n1199), .Z(mult_x_6_n1151) );
  AOI22_X1 U1265 ( .A1(n2185), .A2(n2197), .B1(mul_operand_b_q[15]), .B2(n603), 
        .ZN(n1201) );
  AOI22_X1 U1266 ( .A1(mul_operand_b_q[14]), .A2(n2158), .B1(mult_x_6_n1088), 
        .B2(n1245), .ZN(n1200) );
  NAND2_X1 U1267 ( .A1(n1201), .A2(n1200), .ZN(n1202) );
  XOR2_X1 U1268 ( .A(mul_operand_a_q[29]), .B(n1202), .Z(mult_x_6_n1152) );
  AOI22_X1 U1269 ( .A1(mul_operand_b_q[15]), .A2(n2197), .B1(
        mul_operand_b_q[14]), .B2(n603), .ZN(n1204) );
  AOI22_X1 U1270 ( .A1(mul_operand_b_q[13]), .A2(n2158), .B1(mult_x_6_n1089), 
        .B2(n1245), .ZN(n1203) );
  NAND2_X1 U1271 ( .A1(n1204), .A2(n1203), .ZN(n1205) );
  XOR2_X1 U1272 ( .A(mul_operand_a_q[29]), .B(n1205), .Z(mult_x_6_n1153) );
  AOI22_X1 U1273 ( .A1(mul_operand_b_q[14]), .A2(n2197), .B1(
        mul_operand_b_q[13]), .B2(n603), .ZN(n1207) );
  AOI22_X1 U1274 ( .A1(mul_operand_b_q[12]), .A2(n2158), .B1(n1245), .B2(
        mult_x_6_n1090), .ZN(n1206) );
  NAND2_X1 U1275 ( .A1(n1207), .A2(n1206), .ZN(n1208) );
  XOR2_X1 U1276 ( .A(mul_operand_a_q[29]), .B(n1208), .Z(mult_x_6_n1154) );
  AOI22_X1 U1277 ( .A1(mul_operand_b_q[13]), .A2(n2197), .B1(
        mul_operand_b_q[12]), .B2(n603), .ZN(n1210) );
  AOI22_X1 U1278 ( .A1(mul_operand_b_q[11]), .A2(n2158), .B1(mult_x_6_n1091), 
        .B2(n1245), .ZN(n1209) );
  NAND2_X1 U1279 ( .A1(n1210), .A2(n1209), .ZN(n1211) );
  XOR2_X1 U1280 ( .A(mul_operand_a_q[29]), .B(n1211), .Z(mult_x_6_n1155) );
  AOI22_X1 U1281 ( .A1(mul_operand_b_q[11]), .A2(n603), .B1(
        mul_operand_b_q[12]), .B2(n1246), .ZN(n1213) );
  AOI22_X1 U1282 ( .A1(mul_operand_b_q[10]), .A2(n2158), .B1(mult_x_6_n1092), 
        .B2(n1245), .ZN(n1212) );
  NAND2_X1 U1283 ( .A1(n1213), .A2(n1212), .ZN(n1214) );
  XOR2_X1 U1284 ( .A(mul_operand_a_q[29]), .B(n1214), .Z(mult_x_6_n1156) );
  AOI22_X1 U1285 ( .A1(mul_operand_b_q[11]), .A2(n2197), .B1(
        mul_operand_b_q[10]), .B2(n603), .ZN(n1216) );
  AOI22_X1 U1286 ( .A1(n2187), .A2(n2158), .B1(n2287), .B2(n1245), .ZN(n1215)
         );
  NAND2_X1 U1287 ( .A1(n1216), .A2(n1215), .ZN(n1217) );
  XOR2_X1 U1288 ( .A(mul_operand_a_q[29]), .B(n1217), .Z(mult_x_6_n1157) );
  AOI22_X1 U1289 ( .A1(mul_operand_b_q[10]), .A2(n2197), .B1(n2186), .B2(n603), 
        .ZN(n1219) );
  AOI22_X1 U1290 ( .A1(mul_operand_b_q[8]), .A2(n2158), .B1(mult_x_6_n1094), 
        .B2(n1245), .ZN(n1218) );
  NAND2_X1 U1291 ( .A1(n1219), .A2(n1218), .ZN(n1220) );
  XOR2_X1 U1292 ( .A(mul_operand_a_q[29]), .B(n1220), .Z(mult_x_6_n1158) );
  AOI22_X1 U1293 ( .A1(n2187), .A2(n2197), .B1(mul_operand_b_q[8]), .B2(n603), 
        .ZN(n1222) );
  AOI22_X1 U1294 ( .A1(mul_operand_b_q[7]), .A2(n2158), .B1(mult_x_6_n1095), 
        .B2(n1245), .ZN(n1221) );
  NAND2_X1 U1295 ( .A1(n1222), .A2(n1221), .ZN(n1223) );
  XOR2_X1 U1296 ( .A(mul_operand_a_q[29]), .B(n1223), .Z(mult_x_6_n1159) );
  AOI22_X1 U1297 ( .A1(mul_operand_b_q[8]), .A2(n2197), .B1(mul_operand_b_q[7]), .B2(n603), .ZN(n1225) );
  AOI22_X1 U1298 ( .A1(n2189), .A2(n2158), .B1(n1245), .B2(mult_x_6_n1096), 
        .ZN(n1224) );
  NAND2_X1 U1299 ( .A1(n1225), .A2(n1224), .ZN(n1226) );
  XOR2_X1 U1300 ( .A(mul_operand_a_q[29]), .B(n1226), .Z(mult_x_6_n1160) );
  AOI22_X1 U1301 ( .A1(mul_operand_b_q[7]), .A2(n2197), .B1(n2189), .B2(n603), 
        .ZN(n1228) );
  AOI22_X1 U1302 ( .A1(n2191), .A2(n2158), .B1(n612), .B2(n1245), .ZN(n1227)
         );
  NAND2_X1 U1303 ( .A1(n1228), .A2(n1227), .ZN(n1229) );
  XOR2_X1 U1304 ( .A(mul_operand_a_q[29]), .B(n1229), .Z(mult_x_6_n1161) );
  AOI22_X1 U1305 ( .A1(n2191), .A2(n603), .B1(n2188), .B2(n1246), .ZN(n1231)
         );
  AOI22_X1 U1306 ( .A1(mul_operand_b_q[4]), .A2(n2158), .B1(mult_x_6_n1098), 
        .B2(n1245), .ZN(n1230) );
  NAND2_X1 U1307 ( .A1(n1231), .A2(n1230), .ZN(n1232) );
  XOR2_X1 U1308 ( .A(mul_operand_a_q[29]), .B(n1232), .Z(mult_x_6_n1162) );
  AOI22_X1 U1309 ( .A1(n2191), .A2(n2197), .B1(n2192), .B2(n603), .ZN(n1234)
         );
  AOI22_X1 U1310 ( .A1(n2193), .A2(n2158), .B1(n355), .B2(n1245), .ZN(n1233)
         );
  NAND2_X1 U1311 ( .A1(n1234), .A2(n1233), .ZN(n1235) );
  XOR2_X1 U1312 ( .A(mul_operand_a_q[29]), .B(n1235), .Z(mult_x_6_n1163) );
  AOI22_X1 U1313 ( .A1(mul_operand_b_q[4]), .A2(n2197), .B1(n2193), .B2(n603), 
        .ZN(n1237) );
  AOI22_X1 U1314 ( .A1(mul_operand_b_q[2]), .A2(n2158), .B1(n622), .B2(n1245), 
        .ZN(n1236) );
  NAND2_X1 U1315 ( .A1(n1237), .A2(n1236), .ZN(n1238) );
  XOR2_X1 U1316 ( .A(mul_operand_a_q[29]), .B(n1238), .Z(mult_x_6_n1164) );
  AOI22_X1 U1317 ( .A1(n2193), .A2(n2197), .B1(n1009), .B2(n603), .ZN(n1240)
         );
  AOI22_X1 U1318 ( .A1(n2286), .A2(n2158), .B1(n833), .B2(n1245), .ZN(n1239)
         );
  NAND2_X1 U1319 ( .A1(n1240), .A2(n1239), .ZN(n1241) );
  XOR2_X1 U1320 ( .A(mul_operand_a_q[29]), .B(n1241), .Z(mult_x_6_n1165) );
  AOI22_X1 U1321 ( .A1(n1009), .A2(n2197), .B1(n2195), .B2(n603), .ZN(n1243)
         );
  AOI22_X1 U1322 ( .A1(n1018), .A2(n2158), .B1(mult_x_6_n1102), .B2(n1245), 
        .ZN(n1242) );
  NAND2_X1 U1323 ( .A1(n1243), .A2(n1242), .ZN(n1244) );
  XOR2_X1 U1324 ( .A(mul_operand_a_q[29]), .B(n1244), .Z(mult_x_6_n1166) );
  AOI222_X1 U1325 ( .A1(n2195), .A2(n1246), .B1(n1018), .B2(n603), .C1(n1245), 
        .C2(mult_x_6_n1103), .ZN(n1247) );
  XNOR2_X1 U1326 ( .A(mul_operand_a_q[29]), .B(n1247), .ZN(mult_x_6_n1167) );
  NAND2_X1 U1327 ( .A1(n2157), .A2(n1018), .ZN(n1248) );
  XNOR2_X1 U1328 ( .A(n1248), .B(mul_operand_a_q[29]), .ZN(mult_x_6_n1168) );
  XNOR2_X1 U1329 ( .A(mul_operand_a_q[23]), .B(mul_operand_a_q[24]), .ZN(n1252) );
  XOR2_X1 U1330 ( .A(mul_operand_a_q[26]), .B(mul_operand_a_q[25]), .Z(n1253)
         );
  XNOR2_X1 U1331 ( .A(mul_operand_a_q[25]), .B(mul_operand_a_q[24]), .ZN(n1249) );
  NAND3_X1 U1332 ( .A1(n1253), .A2(n1252), .A3(n1249), .ZN(n1254) );
  NAND3_X1 U1333 ( .A1(n1252), .A2(n1254), .A3(n2417), .ZN(n1250) );
  NAND2_X1 U1334 ( .A1(n1250), .A2(n2177), .ZN(n1251) );
  XOR2_X1 U1335 ( .A(mul_operand_a_q[26]), .B(n1251), .Z(mult_x_6_n1169) );
  NOR2_X1 U1336 ( .A1(n1252), .A2(n1253), .ZN(n1351) );
  OR2_X1 U1337 ( .A1(n1351), .A2(n2198), .ZN(n1255) );
  AOI222_X1 U1338 ( .A1(n1255), .A2(mul_operand_b_q[32]), .B1(mult_x_6_n1071), 
        .B2(n1350), .C1(mul_operand_b_q[31]), .C2(n2156), .ZN(n1256) );
  XNOR2_X1 U1339 ( .A(mul_operand_a_q[26]), .B(n1256), .ZN(mult_x_6_n1170) );
  AOI22_X1 U1340 ( .A1(n2180), .A2(n2156), .B1(mult_x_6_n1072), .B2(n1350), 
        .ZN(n1258) );
  NAND2_X1 U1341 ( .A1(n2177), .A2(n1351), .ZN(n1257) );
  OAI211_X1 U1342 ( .C1(n2178), .C2(n2417), .A(n1258), .B(n1257), .ZN(n1259)
         );
  XOR2_X1 U1343 ( .A(mul_operand_a_q[26]), .B(n1259), .Z(mult_x_6_n1171) );
  AOI22_X1 U1344 ( .A1(n2179), .A2(n1351), .B1(n2180), .B2(n2198), .ZN(n1261)
         );
  AOI22_X1 U1345 ( .A1(mul_operand_b_q[29]), .A2(n2156), .B1(mult_x_6_n1073), 
        .B2(n1350), .ZN(n1260) );
  NAND2_X1 U1346 ( .A1(n1261), .A2(n1260), .ZN(n1262) );
  XOR2_X1 U1347 ( .A(mul_operand_a_q[26]), .B(n1262), .Z(mult_x_6_n1172) );
  AOI22_X1 U1348 ( .A1(n2180), .A2(n1351), .B1(mul_operand_b_q[29]), .B2(n2198), .ZN(n1264) );
  AOI22_X1 U1349 ( .A1(n2181), .A2(n2156), .B1(mult_x_6_n1074), .B2(n1350), 
        .ZN(n1263) );
  NAND2_X1 U1350 ( .A1(n1264), .A2(n1263), .ZN(n1265) );
  XOR2_X1 U1351 ( .A(mul_operand_a_q[26]), .B(n1265), .Z(mult_x_6_n1173) );
  AOI22_X1 U1352 ( .A1(mul_operand_b_q[29]), .A2(n1351), .B1(
        mul_operand_b_q[28]), .B2(n2198), .ZN(n1267) );
  AOI22_X1 U1353 ( .A1(mul_operand_b_q[27]), .A2(n2156), .B1(mult_x_6_n1075), 
        .B2(n1350), .ZN(n1266) );
  NAND2_X1 U1354 ( .A1(n1267), .A2(n1266), .ZN(n1268) );
  XOR2_X1 U1355 ( .A(mul_operand_a_q[26]), .B(n1268), .Z(mult_x_6_n1174) );
  AOI22_X1 U1356 ( .A1(n2181), .A2(n2199), .B1(mul_operand_b_q[27]), .B2(n2198), .ZN(n1270) );
  AOI22_X1 U1357 ( .A1(n2182), .A2(n2156), .B1(mult_x_6_n1076), .B2(n1350), 
        .ZN(n1269) );
  NAND2_X1 U1358 ( .A1(n1270), .A2(n1269), .ZN(n1271) );
  XOR2_X1 U1359 ( .A(mul_operand_a_q[26]), .B(n1271), .Z(mult_x_6_n1175) );
  AOI22_X1 U1360 ( .A1(mul_operand_b_q[27]), .A2(n2199), .B1(
        mul_operand_b_q[26]), .B2(n2198), .ZN(n1273) );
  AOI22_X1 U1361 ( .A1(mul_operand_b_q[25]), .A2(n2156), .B1(mult_x_6_n1077), 
        .B2(n1350), .ZN(n1272) );
  NAND2_X1 U1362 ( .A1(n1273), .A2(n1272), .ZN(n1274) );
  XOR2_X1 U1363 ( .A(mul_operand_a_q[26]), .B(n1274), .Z(mult_x_6_n1176) );
  AOI22_X1 U1364 ( .A1(n2182), .A2(n2199), .B1(mul_operand_b_q[25]), .B2(n2198), .ZN(n1276) );
  AOI22_X1 U1365 ( .A1(n2183), .A2(n2156), .B1(mult_x_6_n1078), .B2(n1350), 
        .ZN(n1275) );
  NAND2_X1 U1366 ( .A1(n1276), .A2(n1275), .ZN(n1277) );
  XOR2_X1 U1367 ( .A(mul_operand_a_q[26]), .B(n1277), .Z(mult_x_6_n1177) );
  AOI22_X1 U1368 ( .A1(mul_operand_b_q[25]), .A2(n2199), .B1(
        mul_operand_b_q[24]), .B2(n626), .ZN(n1279) );
  AOI22_X1 U1369 ( .A1(mul_operand_b_q[23]), .A2(n2156), .B1(mult_x_6_n1079), 
        .B2(n623), .ZN(n1278) );
  NAND2_X1 U1370 ( .A1(n1279), .A2(n1278), .ZN(n1280) );
  XOR2_X1 U1371 ( .A(mul_operand_a_q[26]), .B(n1280), .Z(mult_x_6_n1178) );
  AOI22_X1 U1372 ( .A1(n2183), .A2(n2199), .B1(mul_operand_b_q[23]), .B2(n626), 
        .ZN(n1282) );
  AOI22_X1 U1373 ( .A1(mul_operand_b_q[22]), .A2(n2156), .B1(mult_x_6_n1080), 
        .B2(n623), .ZN(n1281) );
  NAND2_X1 U1374 ( .A1(n1282), .A2(n1281), .ZN(n1283) );
  XOR2_X1 U1375 ( .A(mul_operand_a_q[26]), .B(n1283), .Z(mult_x_6_n1179) );
  AOI22_X1 U1376 ( .A1(mul_operand_b_q[23]), .A2(n2199), .B1(
        mul_operand_b_q[22]), .B2(n626), .ZN(n1285) );
  AOI22_X1 U1377 ( .A1(mul_operand_b_q[21]), .A2(n2156), .B1(mult_x_6_n1081), 
        .B2(n623), .ZN(n1284) );
  NAND2_X1 U1378 ( .A1(n1285), .A2(n1284), .ZN(n1286) );
  XOR2_X1 U1379 ( .A(mul_operand_a_q[26]), .B(n1286), .Z(mult_x_6_n1180) );
  AOI22_X1 U1380 ( .A1(mul_operand_b_q[22]), .A2(n2199), .B1(
        mul_operand_b_q[21]), .B2(n626), .ZN(n1288) );
  AOI22_X1 U1381 ( .A1(mul_operand_b_q[20]), .A2(n2156), .B1(mult_x_6_n1082), 
        .B2(n623), .ZN(n1287) );
  NAND2_X1 U1382 ( .A1(n1288), .A2(n1287), .ZN(n1289) );
  XOR2_X1 U1383 ( .A(mul_operand_a_q[26]), .B(n1289), .Z(mult_x_6_n1181) );
  AOI22_X1 U1384 ( .A1(mul_operand_b_q[21]), .A2(n2199), .B1(
        mul_operand_b_q[20]), .B2(n626), .ZN(n1291) );
  AOI22_X1 U1385 ( .A1(mul_operand_b_q[19]), .A2(n2156), .B1(mult_x_6_n1083), 
        .B2(n623), .ZN(n1290) );
  NAND2_X1 U1386 ( .A1(n1291), .A2(n1290), .ZN(n1292) );
  XOR2_X1 U1387 ( .A(mul_operand_a_q[26]), .B(n1292), .Z(mult_x_6_n1182) );
  AOI22_X1 U1388 ( .A1(mul_operand_b_q[20]), .A2(n2199), .B1(
        mul_operand_b_q[19]), .B2(n626), .ZN(n1294) );
  AOI22_X1 U1389 ( .A1(mul_operand_b_q[18]), .A2(n2156), .B1(mult_x_6_n1084), 
        .B2(n623), .ZN(n1293) );
  NAND2_X1 U1390 ( .A1(n1294), .A2(n1293), .ZN(n1295) );
  XOR2_X1 U1391 ( .A(mul_operand_a_q[26]), .B(n1295), .Z(mult_x_6_n1183) );
  AOI22_X1 U1392 ( .A1(mul_operand_b_q[19]), .A2(n2199), .B1(
        mul_operand_b_q[18]), .B2(n626), .ZN(n1297) );
  AOI22_X1 U1393 ( .A1(mul_operand_b_q[17]), .A2(n2156), .B1(mult_x_6_n1085), 
        .B2(n623), .ZN(n1296) );
  NAND2_X1 U1394 ( .A1(n1297), .A2(n1296), .ZN(n1298) );
  XOR2_X1 U1395 ( .A(mul_operand_a_q[26]), .B(n1298), .Z(mult_x_6_n1184) );
  AOI22_X1 U1396 ( .A1(mul_operand_b_q[17]), .A2(n626), .B1(
        mul_operand_b_q[18]), .B2(n1351), .ZN(n1300) );
  AOI22_X1 U1397 ( .A1(n2185), .A2(n2156), .B1(mult_x_6_n1086), .B2(n623), 
        .ZN(n1299) );
  NAND2_X1 U1398 ( .A1(n1300), .A2(n1299), .ZN(n1301) );
  XOR2_X1 U1399 ( .A(mul_operand_a_q[26]), .B(n1301), .Z(mult_x_6_n1185) );
  AOI22_X1 U1400 ( .A1(mul_operand_b_q[17]), .A2(n2199), .B1(n2184), .B2(n626), 
        .ZN(n1303) );
  AOI22_X1 U1401 ( .A1(mul_operand_b_q[15]), .A2(n2156), .B1(mult_x_6_n1087), 
        .B2(n623), .ZN(n1302) );
  NAND2_X1 U1402 ( .A1(n1303), .A2(n1302), .ZN(n1304) );
  XOR2_X1 U1403 ( .A(mul_operand_a_q[26]), .B(n1304), .Z(mult_x_6_n1186) );
  AOI22_X1 U1404 ( .A1(n2185), .A2(n2199), .B1(mul_operand_b_q[15]), .B2(n626), 
        .ZN(n1306) );
  AOI22_X1 U1405 ( .A1(mul_operand_b_q[14]), .A2(n2156), .B1(mult_x_6_n1088), 
        .B2(n623), .ZN(n1305) );
  NAND2_X1 U1406 ( .A1(n1306), .A2(n1305), .ZN(n1307) );
  XOR2_X1 U1407 ( .A(mul_operand_a_q[26]), .B(n1307), .Z(mult_x_6_n1187) );
  AOI22_X1 U1408 ( .A1(mul_operand_b_q[15]), .A2(n2199), .B1(
        mul_operand_b_q[14]), .B2(n626), .ZN(n1309) );
  AOI22_X1 U1409 ( .A1(mul_operand_b_q[13]), .A2(n2156), .B1(mult_x_6_n1089), 
        .B2(n623), .ZN(n1308) );
  NAND2_X1 U1410 ( .A1(n1309), .A2(n1308), .ZN(n1310) );
  XOR2_X1 U1411 ( .A(mul_operand_a_q[26]), .B(n1310), .Z(mult_x_6_n1188) );
  AOI22_X1 U1412 ( .A1(mul_operand_b_q[14]), .A2(n2199), .B1(
        mul_operand_b_q[13]), .B2(n626), .ZN(n1312) );
  AOI22_X1 U1413 ( .A1(mul_operand_b_q[12]), .A2(n2156), .B1(mult_x_6_n1090), 
        .B2(n623), .ZN(n1311) );
  NAND2_X1 U1414 ( .A1(n1312), .A2(n1311), .ZN(n1313) );
  XOR2_X1 U1415 ( .A(mul_operand_a_q[26]), .B(n1313), .Z(mult_x_6_n1189) );
  AOI22_X1 U1416 ( .A1(mul_operand_b_q[13]), .A2(n2199), .B1(
        mul_operand_b_q[12]), .B2(n626), .ZN(n1315) );
  AOI22_X1 U1417 ( .A1(mul_operand_b_q[11]), .A2(n2156), .B1(mult_x_6_n1091), 
        .B2(n623), .ZN(n1314) );
  NAND2_X1 U1418 ( .A1(n1315), .A2(n1314), .ZN(n1316) );
  XOR2_X1 U1419 ( .A(mul_operand_a_q[26]), .B(n1316), .Z(mult_x_6_n1190) );
  AOI22_X1 U1420 ( .A1(mul_operand_b_q[11]), .A2(n626), .B1(
        mul_operand_b_q[12]), .B2(n1351), .ZN(n1318) );
  AOI22_X1 U1421 ( .A1(mul_operand_b_q[10]), .A2(n2156), .B1(mult_x_6_n1092), 
        .B2(n623), .ZN(n1317) );
  NAND2_X1 U1422 ( .A1(n1318), .A2(n1317), .ZN(n1319) );
  XOR2_X1 U1423 ( .A(mul_operand_a_q[26]), .B(n1319), .Z(mult_x_6_n1191) );
  AOI22_X1 U1424 ( .A1(mul_operand_b_q[11]), .A2(n2199), .B1(
        mul_operand_b_q[10]), .B2(n626), .ZN(n1321) );
  AOI22_X1 U1425 ( .A1(n2187), .A2(n2156), .B1(n2287), .B2(n623), .ZN(n1320)
         );
  NAND2_X1 U1426 ( .A1(n1321), .A2(n1320), .ZN(n1322) );
  XOR2_X1 U1427 ( .A(mul_operand_a_q[26]), .B(n1322), .Z(mult_x_6_n1192) );
  AOI22_X1 U1428 ( .A1(mul_operand_b_q[10]), .A2(n2199), .B1(n2186), .B2(n626), 
        .ZN(n1324) );
  AOI22_X1 U1429 ( .A1(mul_operand_b_q[8]), .A2(n2156), .B1(mult_x_6_n1094), 
        .B2(n623), .ZN(n1323) );
  NAND2_X1 U1430 ( .A1(n1324), .A2(n1323), .ZN(n1325) );
  XOR2_X1 U1431 ( .A(mul_operand_a_q[26]), .B(n1325), .Z(mult_x_6_n1193) );
  AOI22_X1 U1432 ( .A1(n2187), .A2(n2199), .B1(mul_operand_b_q[8]), .B2(n626), 
        .ZN(n1327) );
  AOI22_X1 U1433 ( .A1(mul_operand_b_q[7]), .A2(n2156), .B1(mult_x_6_n1095), 
        .B2(n623), .ZN(n1326) );
  NAND2_X1 U1434 ( .A1(n1327), .A2(n1326), .ZN(n1328) );
  XOR2_X1 U1435 ( .A(mul_operand_a_q[26]), .B(n1328), .Z(mult_x_6_n1194) );
  AOI22_X1 U1436 ( .A1(mul_operand_b_q[8]), .A2(n2199), .B1(mul_operand_b_q[7]), .B2(n626), .ZN(n1330) );
  AOI22_X1 U1437 ( .A1(n2189), .A2(n2156), .B1(mult_x_6_n1096), .B2(n623), 
        .ZN(n1329) );
  NAND2_X1 U1438 ( .A1(n1330), .A2(n1329), .ZN(n1331) );
  XOR2_X1 U1439 ( .A(mul_operand_a_q[26]), .B(n1331), .Z(mult_x_6_n1195) );
  AOI22_X1 U1440 ( .A1(mul_operand_b_q[7]), .A2(n2199), .B1(n2188), .B2(n626), 
        .ZN(n1333) );
  AOI22_X1 U1441 ( .A1(n2191), .A2(n2156), .B1(n612), .B2(n623), .ZN(n1332) );
  NAND2_X1 U1442 ( .A1(n1333), .A2(n1332), .ZN(n1334) );
  XOR2_X1 U1443 ( .A(mul_operand_a_q[26]), .B(n1334), .Z(mult_x_6_n1196) );
  AOI22_X1 U1444 ( .A1(n2191), .A2(n626), .B1(n2188), .B2(n1351), .ZN(n1336)
         );
  AOI22_X1 U1445 ( .A1(mul_operand_b_q[4]), .A2(n2156), .B1(mult_x_6_n1098), 
        .B2(n623), .ZN(n1335) );
  NAND2_X1 U1446 ( .A1(n1336), .A2(n1335), .ZN(n1337) );
  XOR2_X1 U1447 ( .A(mul_operand_a_q[26]), .B(n1337), .Z(mult_x_6_n1197) );
  AOI22_X1 U1448 ( .A1(n2191), .A2(n2199), .B1(n2192), .B2(n626), .ZN(n1339)
         );
  AOI22_X1 U1449 ( .A1(n2193), .A2(n2156), .B1(n355), .B2(n623), .ZN(n1338) );
  NAND2_X1 U1450 ( .A1(n1339), .A2(n1338), .ZN(n1340) );
  XOR2_X1 U1451 ( .A(mul_operand_a_q[26]), .B(n1340), .Z(mult_x_6_n1198) );
  AOI22_X1 U1452 ( .A1(mul_operand_b_q[4]), .A2(n2199), .B1(n2193), .B2(n626), 
        .ZN(n1342) );
  AOI22_X1 U1453 ( .A1(n1009), .A2(n2156), .B1(n622), .B2(n623), .ZN(n1341) );
  NAND2_X1 U1454 ( .A1(n1342), .A2(n1341), .ZN(n1343) );
  XOR2_X1 U1455 ( .A(mul_operand_a_q[26]), .B(n1343), .Z(mult_x_6_n1199) );
  AOI22_X1 U1456 ( .A1(n2193), .A2(n2199), .B1(n1009), .B2(n626), .ZN(n1345)
         );
  AOI22_X1 U1457 ( .A1(n2195), .A2(n2156), .B1(n833), .B2(n623), .ZN(n1344) );
  NAND2_X1 U1458 ( .A1(n1345), .A2(n1344), .ZN(n1346) );
  XOR2_X1 U1459 ( .A(mul_operand_a_q[26]), .B(n1346), .Z(mult_x_6_n1200) );
  AOI22_X1 U1460 ( .A1(n1009), .A2(n2199), .B1(n2195), .B2(n626), .ZN(n1348)
         );
  AOI22_X1 U1461 ( .A1(n1018), .A2(n2156), .B1(mult_x_6_n1102), .B2(n623), 
        .ZN(n1347) );
  NAND2_X1 U1462 ( .A1(n1348), .A2(n1347), .ZN(n1349) );
  XOR2_X1 U1463 ( .A(mul_operand_a_q[26]), .B(n1349), .Z(mult_x_6_n1201) );
  AOI222_X1 U1464 ( .A1(n2286), .A2(n1351), .B1(n1018), .B2(n2198), .C1(n1350), 
        .C2(mult_x_6_n1103), .ZN(n1352) );
  XNOR2_X1 U1465 ( .A(mul_operand_a_q[26]), .B(n1352), .ZN(mult_x_6_n1202) );
  NAND2_X1 U1466 ( .A1(n2155), .A2(n1018), .ZN(n1353) );
  XNOR2_X1 U1467 ( .A(n1353), .B(mul_operand_a_q[26]), .ZN(mult_x_6_n1203) );
  XNOR2_X1 U1468 ( .A(mul_operand_a_q[20]), .B(mul_operand_a_q[21]), .ZN(n1357) );
  XOR2_X1 U1469 ( .A(mul_operand_a_q[23]), .B(mul_operand_a_q[22]), .Z(n1358)
         );
  XNOR2_X1 U1470 ( .A(mul_operand_a_q[22]), .B(mul_operand_a_q[21]), .ZN(n1354) );
  NAND3_X1 U1471 ( .A1(n1358), .A2(n1357), .A3(n1354), .ZN(n1359) );
  NAND3_X1 U1472 ( .A1(n1357), .A2(n1359), .A3(n2418), .ZN(n1355) );
  NAND2_X1 U1473 ( .A1(n1355), .A2(mul_operand_b_q[32]), .ZN(n1356) );
  XOR2_X1 U1474 ( .A(mul_operand_a_q[23]), .B(n1356), .Z(mult_x_6_n1204) );
  NOR2_X1 U1475 ( .A1(n1357), .A2(n1358), .ZN(n1456) );
  OR2_X1 U1476 ( .A1(n607), .A2(n627), .ZN(n1360) );
  AOI222_X1 U1477 ( .A1(n1360), .A2(mul_operand_b_q[32]), .B1(mult_x_6_n1071), 
        .B2(n1455), .C1(mul_operand_b_q[31]), .C2(n2154), .ZN(n1361) );
  XNOR2_X1 U1478 ( .A(mul_operand_a_q[23]), .B(n1361), .ZN(mult_x_6_n1205) );
  AOI22_X1 U1479 ( .A1(n2180), .A2(n2154), .B1(mult_x_6_n1072), .B2(n1455), 
        .ZN(n1363) );
  NAND2_X1 U1480 ( .A1(n2177), .A2(n607), .ZN(n1362) );
  OAI211_X1 U1481 ( .C1(n2178), .C2(n2418), .A(n1363), .B(n1362), .ZN(n1364)
         );
  XOR2_X1 U1482 ( .A(mul_operand_a_q[23]), .B(n1364), .Z(mult_x_6_n1206) );
  AOI22_X1 U1483 ( .A1(n2180), .A2(n627), .B1(mul_operand_b_q[29]), .B2(n2154), 
        .ZN(n1366) );
  AOI22_X1 U1484 ( .A1(n2179), .A2(n607), .B1(mult_x_6_n1073), .B2(n1455), 
        .ZN(n1365) );
  NAND2_X1 U1485 ( .A1(n1366), .A2(n1365), .ZN(n1367) );
  XOR2_X1 U1486 ( .A(mul_operand_a_q[23]), .B(n1367), .Z(mult_x_6_n1207) );
  AOI22_X1 U1487 ( .A1(mul_operand_b_q[29]), .A2(n627), .B1(
        mul_operand_b_q[28]), .B2(n2154), .ZN(n1369) );
  AOI22_X1 U1488 ( .A1(n2180), .A2(n607), .B1(mult_x_6_n1074), .B2(n1455), 
        .ZN(n1368) );
  NAND2_X1 U1489 ( .A1(n1369), .A2(n1368), .ZN(n1370) );
  XOR2_X1 U1490 ( .A(mul_operand_a_q[23]), .B(n1370), .Z(mult_x_6_n1208) );
  AOI22_X1 U1491 ( .A1(n2181), .A2(n2200), .B1(mul_operand_b_q[27]), .B2(n2154), .ZN(n1372) );
  AOI22_X1 U1492 ( .A1(mul_operand_b_q[29]), .A2(n607), .B1(mult_x_6_n1075), 
        .B2(n1455), .ZN(n1371) );
  NAND2_X1 U1493 ( .A1(n1372), .A2(n1371), .ZN(n1373) );
  XOR2_X1 U1494 ( .A(mul_operand_a_q[23]), .B(n1373), .Z(mult_x_6_n1209) );
  AOI22_X1 U1495 ( .A1(mul_operand_b_q[27]), .A2(n627), .B1(
        mul_operand_b_q[26]), .B2(n2154), .ZN(n1375) );
  AOI22_X1 U1496 ( .A1(n2181), .A2(n607), .B1(mult_x_6_n1076), .B2(n1455), 
        .ZN(n1374) );
  NAND2_X1 U1497 ( .A1(n1375), .A2(n1374), .ZN(n1376) );
  XOR2_X1 U1498 ( .A(mul_operand_a_q[23]), .B(n1376), .Z(mult_x_6_n1210) );
  AOI22_X1 U1499 ( .A1(n2182), .A2(n2200), .B1(mul_operand_b_q[25]), .B2(n2154), .ZN(n1378) );
  AOI22_X1 U1500 ( .A1(mul_operand_b_q[27]), .A2(n607), .B1(mult_x_6_n1077), 
        .B2(n1455), .ZN(n1377) );
  NAND2_X1 U1501 ( .A1(n1378), .A2(n1377), .ZN(n1379) );
  XOR2_X1 U1502 ( .A(mul_operand_a_q[23]), .B(n1379), .Z(mult_x_6_n1211) );
  AOI22_X1 U1503 ( .A1(mul_operand_b_q[25]), .A2(n2200), .B1(
        mul_operand_b_q[24]), .B2(n2154), .ZN(n1381) );
  AOI22_X1 U1504 ( .A1(n2182), .A2(n607), .B1(mult_x_6_n1078), .B2(n1455), 
        .ZN(n1380) );
  NAND2_X1 U1505 ( .A1(n1381), .A2(n1380), .ZN(n1382) );
  XOR2_X1 U1506 ( .A(mul_operand_a_q[23]), .B(n1382), .Z(mult_x_6_n1212) );
  AOI22_X1 U1507 ( .A1(n2183), .A2(n2200), .B1(mul_operand_b_q[23]), .B2(n2154), .ZN(n1384) );
  AOI22_X1 U1508 ( .A1(mul_operand_b_q[25]), .A2(n607), .B1(mult_x_6_n1079), 
        .B2(n625), .ZN(n1383) );
  NAND2_X1 U1509 ( .A1(n1384), .A2(n1383), .ZN(n1385) );
  XOR2_X1 U1510 ( .A(mul_operand_a_q[23]), .B(n1385), .Z(mult_x_6_n1213) );
  AOI22_X1 U1511 ( .A1(mul_operand_b_q[23]), .A2(n2200), .B1(
        mul_operand_b_q[22]), .B2(n2154), .ZN(n1387) );
  AOI22_X1 U1512 ( .A1(n2183), .A2(n607), .B1(mult_x_6_n1080), .B2(n625), .ZN(
        n1386) );
  NAND2_X1 U1513 ( .A1(n1387), .A2(n1386), .ZN(n1388) );
  XOR2_X1 U1514 ( .A(mul_operand_a_q[23]), .B(n1388), .Z(mult_x_6_n1214) );
  AOI22_X1 U1515 ( .A1(mul_operand_b_q[22]), .A2(n2200), .B1(
        mul_operand_b_q[21]), .B2(n2154), .ZN(n1390) );
  AOI22_X1 U1516 ( .A1(mul_operand_b_q[23]), .A2(n607), .B1(mult_x_6_n1081), 
        .B2(n625), .ZN(n1389) );
  NAND2_X1 U1517 ( .A1(n1390), .A2(n1389), .ZN(n1391) );
  XOR2_X1 U1518 ( .A(mul_operand_a_q[23]), .B(n1391), .Z(mult_x_6_n1215) );
  AOI22_X1 U1519 ( .A1(mul_operand_b_q[21]), .A2(n2200), .B1(
        mul_operand_b_q[20]), .B2(n2154), .ZN(n1393) );
  AOI22_X1 U1520 ( .A1(mul_operand_b_q[22]), .A2(n607), .B1(mult_x_6_n1082), 
        .B2(n625), .ZN(n1392) );
  NAND2_X1 U1521 ( .A1(n1393), .A2(n1392), .ZN(n1394) );
  XOR2_X1 U1522 ( .A(mul_operand_a_q[23]), .B(n1394), .Z(mult_x_6_n1216) );
  AOI22_X1 U1523 ( .A1(mul_operand_b_q[20]), .A2(n2200), .B1(
        mul_operand_b_q[19]), .B2(n2154), .ZN(n1396) );
  AOI22_X1 U1524 ( .A1(mul_operand_b_q[21]), .A2(n607), .B1(mult_x_6_n1083), 
        .B2(n625), .ZN(n1395) );
  NAND2_X1 U1525 ( .A1(n1396), .A2(n1395), .ZN(n1397) );
  XOR2_X1 U1526 ( .A(mul_operand_a_q[23]), .B(n1397), .Z(mult_x_6_n1217) );
  AOI22_X1 U1527 ( .A1(mul_operand_b_q[19]), .A2(n2200), .B1(
        mul_operand_b_q[18]), .B2(n2154), .ZN(n1399) );
  AOI22_X1 U1528 ( .A1(mul_operand_b_q[20]), .A2(n607), .B1(mult_x_6_n1084), 
        .B2(n625), .ZN(n1398) );
  NAND2_X1 U1529 ( .A1(n1399), .A2(n1398), .ZN(n1400) );
  XOR2_X1 U1530 ( .A(mul_operand_a_q[23]), .B(n1400), .Z(mult_x_6_n1218) );
  AOI22_X1 U1531 ( .A1(mul_operand_b_q[17]), .A2(n2154), .B1(
        mul_operand_b_q[18]), .B2(n627), .ZN(n1402) );
  AOI22_X1 U1532 ( .A1(mul_operand_b_q[19]), .A2(n607), .B1(mult_x_6_n1085), 
        .B2(n625), .ZN(n1401) );
  NAND2_X1 U1533 ( .A1(n1402), .A2(n1401), .ZN(n1403) );
  XOR2_X1 U1534 ( .A(mul_operand_a_q[23]), .B(n1403), .Z(mult_x_6_n1219) );
  AOI22_X1 U1535 ( .A1(mul_operand_b_q[17]), .A2(n2200), .B1(n2184), .B2(n2154), .ZN(n1405) );
  AOI22_X1 U1536 ( .A1(mul_operand_b_q[18]), .A2(n607), .B1(mult_x_6_n1086), 
        .B2(n625), .ZN(n1404) );
  NAND2_X1 U1537 ( .A1(n1405), .A2(n1404), .ZN(n1406) );
  XOR2_X1 U1538 ( .A(mul_operand_a_q[23]), .B(n1406), .Z(mult_x_6_n1220) );
  AOI22_X1 U1539 ( .A1(n2185), .A2(n2200), .B1(mul_operand_b_q[15]), .B2(n2154), .ZN(n1408) );
  AOI22_X1 U1540 ( .A1(mul_operand_b_q[17]), .A2(n607), .B1(mult_x_6_n1087), 
        .B2(n625), .ZN(n1407) );
  NAND2_X1 U1541 ( .A1(n1408), .A2(n1407), .ZN(n1409) );
  XOR2_X1 U1542 ( .A(mul_operand_a_q[23]), .B(n1409), .Z(mult_x_6_n1221) );
  AOI22_X1 U1543 ( .A1(mul_operand_b_q[15]), .A2(n627), .B1(
        mul_operand_b_q[14]), .B2(n2154), .ZN(n1411) );
  AOI22_X1 U1544 ( .A1(n2185), .A2(n607), .B1(mult_x_6_n1088), .B2(n625), .ZN(
        n1410) );
  NAND2_X1 U1545 ( .A1(n1411), .A2(n1410), .ZN(n1412) );
  XOR2_X1 U1546 ( .A(mul_operand_a_q[23]), .B(n1412), .Z(mult_x_6_n1222) );
  AOI22_X1 U1547 ( .A1(mul_operand_b_q[14]), .A2(n627), .B1(
        mul_operand_b_q[13]), .B2(n2154), .ZN(n1414) );
  AOI22_X1 U1548 ( .A1(mul_operand_b_q[15]), .A2(n607), .B1(mult_x_6_n1089), 
        .B2(n625), .ZN(n1413) );
  NAND2_X1 U1549 ( .A1(n1414), .A2(n1413), .ZN(n1415) );
  XOR2_X1 U1550 ( .A(mul_operand_a_q[23]), .B(n1415), .Z(mult_x_6_n1223) );
  AOI22_X1 U1551 ( .A1(mul_operand_b_q[13]), .A2(n627), .B1(
        mul_operand_b_q[12]), .B2(n2154), .ZN(n1417) );
  AOI22_X1 U1552 ( .A1(mul_operand_b_q[14]), .A2(n607), .B1(mult_x_6_n1090), 
        .B2(n625), .ZN(n1416) );
  NAND2_X1 U1553 ( .A1(n1417), .A2(n1416), .ZN(n1418) );
  XOR2_X1 U1554 ( .A(mul_operand_a_q[23]), .B(n1418), .Z(mult_x_6_n1224) );
  AOI22_X1 U1555 ( .A1(mul_operand_b_q[11]), .A2(n2154), .B1(
        mul_operand_b_q[12]), .B2(n627), .ZN(n1420) );
  AOI22_X1 U1556 ( .A1(mul_operand_b_q[13]), .A2(n607), .B1(mult_x_6_n1091), 
        .B2(n625), .ZN(n1419) );
  NAND2_X1 U1557 ( .A1(n1420), .A2(n1419), .ZN(n1421) );
  XOR2_X1 U1558 ( .A(mul_operand_a_q[23]), .B(n1421), .Z(mult_x_6_n1225) );
  AOI22_X1 U1559 ( .A1(mul_operand_b_q[11]), .A2(n627), .B1(
        mul_operand_b_q[10]), .B2(n2154), .ZN(n1423) );
  AOI22_X1 U1560 ( .A1(mul_operand_b_q[12]), .A2(n607), .B1(mult_x_6_n1092), 
        .B2(n625), .ZN(n1422) );
  NAND2_X1 U1561 ( .A1(n1423), .A2(n1422), .ZN(n1424) );
  XOR2_X1 U1562 ( .A(mul_operand_a_q[23]), .B(n1424), .Z(mult_x_6_n1226) );
  AOI22_X1 U1563 ( .A1(mul_operand_b_q[10]), .A2(n627), .B1(n2186), .B2(n2154), 
        .ZN(n1426) );
  AOI22_X1 U1564 ( .A1(mul_operand_b_q[11]), .A2(n607), .B1(n2287), .B2(n625), 
        .ZN(n1425) );
  NAND2_X1 U1565 ( .A1(n1426), .A2(n1425), .ZN(n1427) );
  XOR2_X1 U1566 ( .A(mul_operand_a_q[23]), .B(n1427), .Z(mult_x_6_n1227) );
  AOI22_X1 U1567 ( .A1(n2187), .A2(n627), .B1(mul_operand_b_q[8]), .B2(n2154), 
        .ZN(n1429) );
  AOI22_X1 U1568 ( .A1(mul_operand_b_q[10]), .A2(n607), .B1(mult_x_6_n1094), 
        .B2(n625), .ZN(n1428) );
  NAND2_X1 U1569 ( .A1(n1429), .A2(n1428), .ZN(n1430) );
  XOR2_X1 U1570 ( .A(mul_operand_a_q[23]), .B(n1430), .Z(mult_x_6_n1228) );
  AOI22_X1 U1571 ( .A1(mul_operand_b_q[8]), .A2(n2200), .B1(mul_operand_b_q[7]), .B2(n2154), .ZN(n1432) );
  AOI22_X1 U1572 ( .A1(n2187), .A2(n607), .B1(mult_x_6_n1095), .B2(n625), .ZN(
        n1431) );
  NAND2_X1 U1573 ( .A1(n1432), .A2(n1431), .ZN(n1433) );
  XOR2_X1 U1574 ( .A(mul_operand_a_q[23]), .B(n1433), .Z(mult_x_6_n1229) );
  AOI22_X1 U1575 ( .A1(mul_operand_b_q[7]), .A2(n627), .B1(n2188), .B2(n2154), 
        .ZN(n1435) );
  AOI22_X1 U1576 ( .A1(mul_operand_b_q[8]), .A2(n607), .B1(mult_x_6_n1096), 
        .B2(n625), .ZN(n1434) );
  NAND2_X1 U1577 ( .A1(n1435), .A2(n1434), .ZN(n1436) );
  XOR2_X1 U1578 ( .A(mul_operand_a_q[23]), .B(n1436), .Z(mult_x_6_n1230) );
  AOI22_X1 U1579 ( .A1(n2191), .A2(n2154), .B1(n2188), .B2(n627), .ZN(n1438)
         );
  AOI22_X1 U1580 ( .A1(mul_operand_b_q[7]), .A2(n607), .B1(n612), .B2(n625), 
        .ZN(n1437) );
  NAND2_X1 U1581 ( .A1(n1438), .A2(n1437), .ZN(n1439) );
  XOR2_X1 U1582 ( .A(mul_operand_a_q[23]), .B(n1439), .Z(mult_x_6_n1231) );
  AOI22_X1 U1583 ( .A1(n2191), .A2(n627), .B1(n2192), .B2(n2154), .ZN(n1441)
         );
  AOI22_X1 U1584 ( .A1(n2189), .A2(n607), .B1(mult_x_6_n1098), .B2(n625), .ZN(
        n1440) );
  NAND2_X1 U1585 ( .A1(n1441), .A2(n1440), .ZN(n1442) );
  XOR2_X1 U1586 ( .A(mul_operand_a_q[23]), .B(n1442), .Z(mult_x_6_n1232) );
  AOI22_X1 U1587 ( .A1(mul_operand_b_q[4]), .A2(n627), .B1(n2193), .B2(n2154), 
        .ZN(n1444) );
  AOI22_X1 U1588 ( .A1(n2191), .A2(n607), .B1(n355), .B2(n625), .ZN(n1443) );
  NAND2_X1 U1589 ( .A1(n1444), .A2(n1443), .ZN(n1445) );
  XOR2_X1 U1590 ( .A(mul_operand_a_q[23]), .B(n1445), .Z(mult_x_6_n1233) );
  AOI22_X1 U1591 ( .A1(n2193), .A2(n627), .B1(n1009), .B2(n2154), .ZN(n1447)
         );
  AOI22_X1 U1592 ( .A1(mul_operand_b_q[4]), .A2(n607), .B1(n622), .B2(n625), 
        .ZN(n1446) );
  NAND2_X1 U1593 ( .A1(n1447), .A2(n1446), .ZN(n1448) );
  XOR2_X1 U1594 ( .A(mul_operand_a_q[23]), .B(n1448), .Z(mult_x_6_n1234) );
  AOI22_X1 U1595 ( .A1(mul_operand_b_q[2]), .A2(n627), .B1(n2195), .B2(n2154), 
        .ZN(n1450) );
  AOI22_X1 U1596 ( .A1(n2193), .A2(n607), .B1(n833), .B2(n625), .ZN(n1449) );
  NAND2_X1 U1597 ( .A1(n1450), .A2(n1449), .ZN(n1451) );
  XOR2_X1 U1598 ( .A(mul_operand_a_q[23]), .B(n1451), .Z(mult_x_6_n1235) );
  AOI22_X1 U1599 ( .A1(n2195), .A2(n627), .B1(n1018), .B2(n2154), .ZN(n1453)
         );
  AOI22_X1 U1600 ( .A1(n1009), .A2(n607), .B1(mult_x_6_n1102), .B2(n625), .ZN(
        n1452) );
  NAND2_X1 U1601 ( .A1(n1453), .A2(n1452), .ZN(n1454) );
  XOR2_X1 U1602 ( .A(mul_operand_a_q[23]), .B(n1454), .Z(mult_x_6_n1236) );
  AOI222_X1 U1603 ( .A1(n2286), .A2(n1456), .B1(n1018), .B2(n627), .C1(n1455), 
        .C2(mult_x_6_n1103), .ZN(n1457) );
  XNOR2_X1 U1604 ( .A(mul_operand_a_q[23]), .B(n1457), .ZN(mult_x_6_n1237) );
  NAND2_X1 U1605 ( .A1(n2153), .A2(n1018), .ZN(n1458) );
  XNOR2_X1 U1606 ( .A(n1458), .B(mul_operand_a_q[23]), .ZN(mult_x_6_n1238) );
  XNOR2_X1 U1607 ( .A(mul_operand_a_q[17]), .B(mul_operand_a_q[18]), .ZN(n1462) );
  XOR2_X1 U1608 ( .A(mul_operand_a_q[20]), .B(mul_operand_a_q[19]), .Z(n1463)
         );
  XNOR2_X1 U1609 ( .A(mul_operand_a_q[19]), .B(mul_operand_a_q[18]), .ZN(n1459) );
  NAND3_X1 U1610 ( .A1(n1463), .A2(n1462), .A3(n1459), .ZN(n1464) );
  NAND3_X1 U1611 ( .A1(n1462), .A2(n1464), .A3(n2419), .ZN(n1460) );
  NAND2_X1 U1612 ( .A1(n1460), .A2(mul_operand_b_q[32]), .ZN(n1461) );
  XOR2_X1 U1613 ( .A(n2170), .B(n1461), .Z(mult_x_6_n1239) );
  NOR2_X1 U1614 ( .A1(n1462), .A2(n1463), .ZN(n1561) );
  OR2_X1 U1615 ( .A1(n1561), .A2(n2202), .ZN(n1465) );
  AOI222_X1 U1616 ( .A1(n1465), .A2(mul_operand_b_q[32]), .B1(mult_x_6_n1071), 
        .B2(n1560), .C1(n2179), .C2(n2152), .ZN(n1466) );
  XNOR2_X1 U1617 ( .A(n2170), .B(n1466), .ZN(mult_x_6_n1240) );
  AOI22_X1 U1618 ( .A1(n2180), .A2(n2152), .B1(mult_x_6_n1072), .B2(n1560), 
        .ZN(n1468) );
  NAND2_X1 U1619 ( .A1(n2177), .A2(n1561), .ZN(n1467) );
  OAI211_X1 U1620 ( .C1(n2178), .C2(n2419), .A(n1468), .B(n1467), .ZN(n1469)
         );
  XOR2_X1 U1621 ( .A(n2170), .B(n1469), .Z(mult_x_6_n1241) );
  AOI22_X1 U1622 ( .A1(n2179), .A2(n1561), .B1(n2180), .B2(n2202), .ZN(n1471)
         );
  AOI22_X1 U1623 ( .A1(mul_operand_b_q[29]), .A2(n2152), .B1(mult_x_6_n1073), 
        .B2(n1560), .ZN(n1470) );
  NAND2_X1 U1624 ( .A1(n1471), .A2(n1470), .ZN(n1472) );
  XOR2_X1 U1625 ( .A(n2170), .B(n1472), .Z(mult_x_6_n1242) );
  AOI22_X1 U1626 ( .A1(n2180), .A2(n1561), .B1(mul_operand_b_q[29]), .B2(n2202), .ZN(n1474) );
  AOI22_X1 U1627 ( .A1(n2181), .A2(n2152), .B1(mult_x_6_n1074), .B2(n1560), 
        .ZN(n1473) );
  NAND2_X1 U1628 ( .A1(n1474), .A2(n1473), .ZN(n1475) );
  XOR2_X1 U1629 ( .A(n2170), .B(n1475), .Z(mult_x_6_n1243) );
  AOI22_X1 U1630 ( .A1(mul_operand_b_q[29]), .A2(n1561), .B1(
        mul_operand_b_q[28]), .B2(n2202), .ZN(n1477) );
  AOI22_X1 U1631 ( .A1(mul_operand_b_q[27]), .A2(n2152), .B1(mult_x_6_n1075), 
        .B2(n1560), .ZN(n1476) );
  NAND2_X1 U1632 ( .A1(n1477), .A2(n1476), .ZN(n1478) );
  XOR2_X1 U1633 ( .A(n2170), .B(n1478), .Z(mult_x_6_n1244) );
  AOI22_X1 U1634 ( .A1(n2181), .A2(n631), .B1(mul_operand_b_q[27]), .B2(n2202), 
        .ZN(n1480) );
  AOI22_X1 U1635 ( .A1(n2182), .A2(n2152), .B1(mult_x_6_n1076), .B2(n1560), 
        .ZN(n1479) );
  NAND2_X1 U1636 ( .A1(n1480), .A2(n1479), .ZN(n1481) );
  XOR2_X1 U1637 ( .A(n2170), .B(n1481), .Z(mult_x_6_n1245) );
  AOI22_X1 U1638 ( .A1(mul_operand_b_q[27]), .A2(n631), .B1(
        mul_operand_b_q[26]), .B2(n2202), .ZN(n1483) );
  AOI22_X1 U1639 ( .A1(mul_operand_b_q[25]), .A2(n2152), .B1(mult_x_6_n1077), 
        .B2(n1560), .ZN(n1482) );
  NAND2_X1 U1640 ( .A1(n1483), .A2(n1482), .ZN(n1484) );
  XOR2_X1 U1641 ( .A(n2170), .B(n1484), .Z(mult_x_6_n1246) );
  AOI22_X1 U1642 ( .A1(n2182), .A2(n631), .B1(mul_operand_b_q[25]), .B2(n2202), 
        .ZN(n1486) );
  AOI22_X1 U1643 ( .A1(n2183), .A2(n2152), .B1(mult_x_6_n1078), .B2(n1560), 
        .ZN(n1485) );
  NAND2_X1 U1644 ( .A1(n1486), .A2(n1485), .ZN(n1487) );
  XOR2_X1 U1645 ( .A(n2170), .B(n1487), .Z(mult_x_6_n1247) );
  AOI22_X1 U1646 ( .A1(mul_operand_b_q[25]), .A2(n631), .B1(
        mul_operand_b_q[24]), .B2(n605), .ZN(n1489) );
  AOI22_X1 U1647 ( .A1(mul_operand_b_q[23]), .A2(n2152), .B1(mult_x_6_n1079), 
        .B2(n2201), .ZN(n1488) );
  NAND2_X1 U1648 ( .A1(n1489), .A2(n1488), .ZN(n1490) );
  XOR2_X1 U1649 ( .A(n2170), .B(n1490), .Z(mult_x_6_n1248) );
  AOI22_X1 U1650 ( .A1(n2183), .A2(n631), .B1(mul_operand_b_q[23]), .B2(n605), 
        .ZN(n1492) );
  AOI22_X1 U1651 ( .A1(mul_operand_b_q[22]), .A2(n2152), .B1(mult_x_6_n1080), 
        .B2(n2201), .ZN(n1491) );
  NAND2_X1 U1652 ( .A1(n1492), .A2(n1491), .ZN(n1493) );
  XOR2_X1 U1653 ( .A(n2170), .B(n1493), .Z(mult_x_6_n1249) );
  AOI22_X1 U1654 ( .A1(mul_operand_b_q[23]), .A2(n631), .B1(
        mul_operand_b_q[22]), .B2(n605), .ZN(n1495) );
  AOI22_X1 U1655 ( .A1(mul_operand_b_q[21]), .A2(n2152), .B1(mult_x_6_n1081), 
        .B2(n2201), .ZN(n1494) );
  NAND2_X1 U1656 ( .A1(n1495), .A2(n1494), .ZN(n1496) );
  XOR2_X1 U1657 ( .A(n2170), .B(n1496), .Z(mult_x_6_n1250) );
  AOI22_X1 U1658 ( .A1(mul_operand_b_q[22]), .A2(n631), .B1(
        mul_operand_b_q[21]), .B2(n605), .ZN(n1498) );
  AOI22_X1 U1659 ( .A1(mul_operand_b_q[20]), .A2(n2152), .B1(mult_x_6_n1082), 
        .B2(n2201), .ZN(n1497) );
  NAND2_X1 U1660 ( .A1(n1498), .A2(n1497), .ZN(n1499) );
  XOR2_X1 U1661 ( .A(n2170), .B(n1499), .Z(mult_x_6_n1251) );
  AOI22_X1 U1662 ( .A1(mul_operand_b_q[21]), .A2(n631), .B1(
        mul_operand_b_q[20]), .B2(n605), .ZN(n1501) );
  AOI22_X1 U1663 ( .A1(mul_operand_b_q[19]), .A2(n2152), .B1(mult_x_6_n1083), 
        .B2(n2201), .ZN(n1500) );
  NAND2_X1 U1664 ( .A1(n1501), .A2(n1500), .ZN(n1502) );
  XOR2_X1 U1665 ( .A(n2170), .B(n1502), .Z(mult_x_6_n1252) );
  AOI22_X1 U1666 ( .A1(mul_operand_b_q[20]), .A2(n631), .B1(
        mul_operand_b_q[19]), .B2(n605), .ZN(n1504) );
  AOI22_X1 U1667 ( .A1(mul_operand_b_q[18]), .A2(n2152), .B1(mult_x_6_n1084), 
        .B2(n2201), .ZN(n1503) );
  NAND2_X1 U1668 ( .A1(n1504), .A2(n1503), .ZN(n1505) );
  XOR2_X1 U1669 ( .A(n2170), .B(n1505), .Z(mult_x_6_n1253) );
  AOI22_X1 U1670 ( .A1(mul_operand_b_q[19]), .A2(n631), .B1(
        mul_operand_b_q[18]), .B2(n605), .ZN(n1507) );
  AOI22_X1 U1671 ( .A1(mul_operand_b_q[17]), .A2(n2152), .B1(mult_x_6_n1085), 
        .B2(n2201), .ZN(n1506) );
  NAND2_X1 U1672 ( .A1(n1507), .A2(n1506), .ZN(n1508) );
  XOR2_X1 U1673 ( .A(n2170), .B(n1508), .Z(mult_x_6_n1254) );
  AOI22_X1 U1674 ( .A1(mul_operand_b_q[17]), .A2(n605), .B1(
        mul_operand_b_q[18]), .B2(n1561), .ZN(n1510) );
  AOI22_X1 U1675 ( .A1(n2185), .A2(n2152), .B1(mult_x_6_n1086), .B2(n2201), 
        .ZN(n1509) );
  NAND2_X1 U1676 ( .A1(n1510), .A2(n1509), .ZN(n1511) );
  XOR2_X1 U1677 ( .A(n2170), .B(n1511), .Z(mult_x_6_n1255) );
  AOI22_X1 U1678 ( .A1(mul_operand_b_q[17]), .A2(n631), .B1(n2184), .B2(n605), 
        .ZN(n1513) );
  AOI22_X1 U1679 ( .A1(mul_operand_b_q[15]), .A2(n2152), .B1(mult_x_6_n1087), 
        .B2(n2201), .ZN(n1512) );
  NAND2_X1 U1680 ( .A1(n1513), .A2(n1512), .ZN(n1514) );
  XOR2_X1 U1681 ( .A(n2170), .B(n1514), .Z(mult_x_6_n1256) );
  AOI22_X1 U1682 ( .A1(n2185), .A2(n631), .B1(mul_operand_b_q[15]), .B2(n605), 
        .ZN(n1516) );
  AOI22_X1 U1683 ( .A1(mul_operand_b_q[14]), .A2(n2152), .B1(mult_x_6_n1088), 
        .B2(n2201), .ZN(n1515) );
  NAND2_X1 U1684 ( .A1(n1516), .A2(n1515), .ZN(n1517) );
  XOR2_X1 U1685 ( .A(n2170), .B(n1517), .Z(mult_x_6_n1257) );
  AOI22_X1 U1686 ( .A1(mul_operand_b_q[15]), .A2(n631), .B1(
        mul_operand_b_q[14]), .B2(n605), .ZN(n1519) );
  AOI22_X1 U1687 ( .A1(mul_operand_b_q[13]), .A2(n2152), .B1(mult_x_6_n1089), 
        .B2(n2201), .ZN(n1518) );
  NAND2_X1 U1688 ( .A1(n1519), .A2(n1518), .ZN(n1520) );
  XOR2_X1 U1689 ( .A(n2170), .B(n1520), .Z(mult_x_6_n1258) );
  AOI22_X1 U1690 ( .A1(mul_operand_b_q[14]), .A2(n631), .B1(
        mul_operand_b_q[13]), .B2(n605), .ZN(n1522) );
  AOI22_X1 U1691 ( .A1(mul_operand_b_q[12]), .A2(n2152), .B1(mult_x_6_n1090), 
        .B2(n1560), .ZN(n1521) );
  NAND2_X1 U1692 ( .A1(n1522), .A2(n1521), .ZN(n1523) );
  XOR2_X1 U1693 ( .A(n2170), .B(n1523), .Z(mult_x_6_n1259) );
  AOI22_X1 U1694 ( .A1(mul_operand_b_q[13]), .A2(n631), .B1(
        mul_operand_b_q[12]), .B2(n605), .ZN(n1525) );
  AOI22_X1 U1695 ( .A1(mul_operand_b_q[11]), .A2(n2152), .B1(mult_x_6_n1091), 
        .B2(n1560), .ZN(n1524) );
  NAND2_X1 U1696 ( .A1(n1525), .A2(n1524), .ZN(n1526) );
  XOR2_X1 U1697 ( .A(n2170), .B(n1526), .Z(mult_x_6_n1260) );
  AOI22_X1 U1698 ( .A1(mul_operand_b_q[11]), .A2(n605), .B1(
        mul_operand_b_q[12]), .B2(n1561), .ZN(n1528) );
  AOI22_X1 U1699 ( .A1(mul_operand_b_q[10]), .A2(n2152), .B1(mult_x_6_n1092), 
        .B2(n1560), .ZN(n1527) );
  NAND2_X1 U1700 ( .A1(n1528), .A2(n1527), .ZN(n1529) );
  XOR2_X1 U1701 ( .A(n2170), .B(n1529), .Z(mult_x_6_n1261) );
  AOI22_X1 U1702 ( .A1(mul_operand_b_q[11]), .A2(n631), .B1(
        mul_operand_b_q[10]), .B2(n605), .ZN(n1531) );
  AOI22_X1 U1703 ( .A1(n2187), .A2(n2152), .B1(n2287), .B2(n1560), .ZN(n1530)
         );
  NAND2_X1 U1704 ( .A1(n1531), .A2(n1530), .ZN(n1532) );
  XOR2_X1 U1705 ( .A(n2170), .B(n1532), .Z(mult_x_6_n1262) );
  AOI22_X1 U1706 ( .A1(mul_operand_b_q[10]), .A2(n631), .B1(n2186), .B2(n605), 
        .ZN(n1534) );
  AOI22_X1 U1707 ( .A1(mul_operand_b_q[8]), .A2(n2152), .B1(mult_x_6_n1094), 
        .B2(n1560), .ZN(n1533) );
  NAND2_X1 U1708 ( .A1(n1534), .A2(n1533), .ZN(n1535) );
  XOR2_X1 U1709 ( .A(n2170), .B(n1535), .Z(mult_x_6_n1263) );
  AOI22_X1 U1710 ( .A1(n2187), .A2(n631), .B1(mul_operand_b_q[8]), .B2(n605), 
        .ZN(n1537) );
  AOI22_X1 U1711 ( .A1(mul_operand_b_q[7]), .A2(n2152), .B1(mult_x_6_n1095), 
        .B2(n2201), .ZN(n1536) );
  NAND2_X1 U1712 ( .A1(n1537), .A2(n1536), .ZN(n1538) );
  XOR2_X1 U1713 ( .A(n2170), .B(n1538), .Z(mult_x_6_n1264) );
  AOI22_X1 U1714 ( .A1(mul_operand_b_q[8]), .A2(n631), .B1(mul_operand_b_q[7]), 
        .B2(n605), .ZN(n1540) );
  AOI22_X1 U1715 ( .A1(n2189), .A2(n2152), .B1(mult_x_6_n1096), .B2(n1560), 
        .ZN(n1539) );
  NAND2_X1 U1716 ( .A1(n1540), .A2(n1539), .ZN(n1541) );
  XOR2_X1 U1717 ( .A(n2170), .B(n1541), .Z(mult_x_6_n1265) );
  AOI22_X1 U1718 ( .A1(mul_operand_b_q[7]), .A2(n631), .B1(n2188), .B2(n605), 
        .ZN(n1543) );
  AOI22_X1 U1719 ( .A1(n2191), .A2(n2152), .B1(n612), .B2(n1560), .ZN(n1542)
         );
  NAND2_X1 U1720 ( .A1(n1543), .A2(n1542), .ZN(n1544) );
  XOR2_X1 U1721 ( .A(n2170), .B(n1544), .Z(mult_x_6_n1266) );
  AOI22_X1 U1722 ( .A1(n2191), .A2(n605), .B1(n2188), .B2(n1561), .ZN(n1546)
         );
  AOI22_X1 U1723 ( .A1(mul_operand_b_q[4]), .A2(n2152), .B1(mult_x_6_n1098), 
        .B2(n1560), .ZN(n1545) );
  NAND2_X1 U1724 ( .A1(n1546), .A2(n1545), .ZN(n1547) );
  XOR2_X1 U1725 ( .A(n2170), .B(n1547), .Z(mult_x_6_n1267) );
  AOI22_X1 U1726 ( .A1(n2191), .A2(n631), .B1(n2192), .B2(n605), .ZN(n1549) );
  AOI22_X1 U1727 ( .A1(n2193), .A2(n2152), .B1(n355), .B2(n1560), .ZN(n1548)
         );
  NAND2_X1 U1728 ( .A1(n1549), .A2(n1548), .ZN(n1550) );
  XOR2_X1 U1729 ( .A(n2170), .B(n1550), .Z(mult_x_6_n1268) );
  AOI22_X1 U1730 ( .A1(mul_operand_b_q[4]), .A2(n631), .B1(n2193), .B2(n605), 
        .ZN(n1552) );
  AOI22_X1 U1731 ( .A1(n1009), .A2(n2152), .B1(n622), .B2(n1560), .ZN(n1551)
         );
  NAND2_X1 U1732 ( .A1(n1552), .A2(n1551), .ZN(n1553) );
  XOR2_X1 U1733 ( .A(n2170), .B(n1553), .Z(mult_x_6_n1269) );
  AOI22_X1 U1734 ( .A1(n2193), .A2(n631), .B1(n1009), .B2(n605), .ZN(n1555) );
  AOI22_X1 U1735 ( .A1(n2195), .A2(n2152), .B1(n833), .B2(n1560), .ZN(n1554)
         );
  NAND2_X1 U1736 ( .A1(n1555), .A2(n1554), .ZN(n1556) );
  XOR2_X1 U1737 ( .A(n2170), .B(n1556), .Z(mult_x_6_n1270) );
  AOI22_X1 U1738 ( .A1(mul_operand_b_q[2]), .A2(n631), .B1(n2286), .B2(n605), 
        .ZN(n1558) );
  AOI22_X1 U1739 ( .A1(n1018), .A2(n2152), .B1(mult_x_6_n1102), .B2(n1560), 
        .ZN(n1557) );
  NAND2_X1 U1740 ( .A1(n1558), .A2(n1557), .ZN(n1559) );
  XOR2_X1 U1741 ( .A(n2170), .B(n1559), .Z(mult_x_6_n1271) );
  AOI222_X1 U1742 ( .A1(n2195), .A2(n1561), .B1(n1018), .B2(n2202), .C1(n1560), 
        .C2(mult_x_6_n1103), .ZN(n1562) );
  XNOR2_X1 U1743 ( .A(n2170), .B(n1562), .ZN(mult_x_6_n1272) );
  NAND2_X1 U1744 ( .A1(n2151), .A2(n1018), .ZN(n1563) );
  XNOR2_X1 U1745 ( .A(n1563), .B(n2170), .ZN(mult_x_6_n1273) );
  XNOR2_X1 U1746 ( .A(mul_operand_a_q[14]), .B(mul_operand_a_q[15]), .ZN(n1567) );
  XOR2_X1 U1747 ( .A(mul_operand_a_q[17]), .B(mul_operand_a_q[16]), .Z(n1568)
         );
  XNOR2_X1 U1748 ( .A(mul_operand_a_q[16]), .B(mul_operand_a_q[15]), .ZN(n1564) );
  NAND3_X1 U1749 ( .A1(n1568), .A2(n1567), .A3(n1564), .ZN(n1569) );
  NAND3_X1 U1750 ( .A1(n1567), .A2(n1569), .A3(n2425), .ZN(n1565) );
  NAND2_X1 U1751 ( .A1(n1565), .A2(mul_operand_b_q[32]), .ZN(n1566) );
  XOR2_X1 U1752 ( .A(n2171), .B(n1566), .Z(mult_x_6_n1274) );
  NOR2_X1 U1753 ( .A1(n1567), .A2(n1568), .ZN(n1666) );
  OR2_X1 U1754 ( .A1(n1666), .A2(n2203), .ZN(n1570) );
  AOI222_X1 U1755 ( .A1(n1570), .A2(mul_operand_b_q[32]), .B1(mult_x_6_n1071), 
        .B2(n1665), .C1(n2179), .C2(n2150), .ZN(n1571) );
  XNOR2_X1 U1756 ( .A(n2171), .B(n1571), .ZN(mult_x_6_n1275) );
  AOI22_X1 U1757 ( .A1(n2180), .A2(n2150), .B1(mult_x_6_n1072), .B2(n1665), 
        .ZN(n1573) );
  NAND2_X1 U1758 ( .A1(n2177), .A2(n1666), .ZN(n1572) );
  OAI211_X1 U1759 ( .C1(n2178), .C2(n2425), .A(n1573), .B(n1572), .ZN(n1574)
         );
  XOR2_X1 U1760 ( .A(n2171), .B(n1574), .Z(mult_x_6_n1276) );
  AOI22_X1 U1761 ( .A1(n2179), .A2(n1666), .B1(n2180), .B2(n2203), .ZN(n1576)
         );
  AOI22_X1 U1762 ( .A1(mul_operand_b_q[29]), .A2(n2150), .B1(mult_x_6_n1073), 
        .B2(n1665), .ZN(n1575) );
  NAND2_X1 U1763 ( .A1(n1576), .A2(n1575), .ZN(n1577) );
  XOR2_X1 U1764 ( .A(n2171), .B(n1577), .Z(mult_x_6_n1277) );
  AOI22_X1 U1765 ( .A1(n2180), .A2(n1666), .B1(mul_operand_b_q[29]), .B2(n2203), .ZN(n1579) );
  AOI22_X1 U1766 ( .A1(n2181), .A2(n2150), .B1(mult_x_6_n1074), .B2(n1665), 
        .ZN(n1578) );
  NAND2_X1 U1767 ( .A1(n1579), .A2(n1578), .ZN(n1580) );
  XOR2_X1 U1768 ( .A(n2171), .B(n1580), .Z(mult_x_6_n1278) );
  AOI22_X1 U1769 ( .A1(mul_operand_b_q[29]), .A2(n1666), .B1(
        mul_operand_b_q[28]), .B2(n2203), .ZN(n1582) );
  AOI22_X1 U1770 ( .A1(mul_operand_b_q[27]), .A2(n2150), .B1(mult_x_6_n1075), 
        .B2(n1665), .ZN(n1581) );
  NAND2_X1 U1771 ( .A1(n1582), .A2(n1581), .ZN(n1583) );
  XOR2_X1 U1772 ( .A(n2171), .B(n1583), .Z(mult_x_6_n1279) );
  AOI22_X1 U1773 ( .A1(n2181), .A2(n628), .B1(mul_operand_b_q[27]), .B2(n2203), 
        .ZN(n1585) );
  AOI22_X1 U1774 ( .A1(n2182), .A2(n2150), .B1(mult_x_6_n1076), .B2(n1665), 
        .ZN(n1584) );
  NAND2_X1 U1775 ( .A1(n1585), .A2(n1584), .ZN(n1586) );
  XOR2_X1 U1776 ( .A(n2171), .B(n1586), .Z(mult_x_6_n1280) );
  AOI22_X1 U1777 ( .A1(mul_operand_b_q[27]), .A2(n628), .B1(
        mul_operand_b_q[26]), .B2(n2203), .ZN(n1588) );
  AOI22_X1 U1778 ( .A1(mul_operand_b_q[25]), .A2(n2150), .B1(mult_x_6_n1077), 
        .B2(n1665), .ZN(n1587) );
  NAND2_X1 U1779 ( .A1(n1588), .A2(n1587), .ZN(n1589) );
  XOR2_X1 U1780 ( .A(n2171), .B(n1589), .Z(mult_x_6_n1281) );
  AOI22_X1 U1781 ( .A1(n2182), .A2(n628), .B1(mul_operand_b_q[25]), .B2(n2203), 
        .ZN(n1591) );
  AOI22_X1 U1782 ( .A1(n2183), .A2(n2150), .B1(mult_x_6_n1078), .B2(n1665), 
        .ZN(n1590) );
  NAND2_X1 U1783 ( .A1(n1591), .A2(n1590), .ZN(n1592) );
  XOR2_X1 U1784 ( .A(n2171), .B(n1592), .Z(mult_x_6_n1282) );
  AOI22_X1 U1785 ( .A1(mul_operand_b_q[25]), .A2(n628), .B1(
        mul_operand_b_q[24]), .B2(n606), .ZN(n1594) );
  AOI22_X1 U1786 ( .A1(mul_operand_b_q[23]), .A2(n2150), .B1(mult_x_6_n1079), 
        .B2(n1665), .ZN(n1593) );
  NAND2_X1 U1787 ( .A1(n1594), .A2(n1593), .ZN(n1595) );
  XOR2_X1 U1788 ( .A(n2171), .B(n1595), .Z(mult_x_6_n1283) );
  AOI22_X1 U1789 ( .A1(n2183), .A2(n628), .B1(mul_operand_b_q[23]), .B2(n606), 
        .ZN(n1597) );
  AOI22_X1 U1790 ( .A1(mul_operand_b_q[22]), .A2(n2150), .B1(mult_x_6_n1080), 
        .B2(n1665), .ZN(n1596) );
  NAND2_X1 U1791 ( .A1(n1597), .A2(n1596), .ZN(n1598) );
  XOR2_X1 U1792 ( .A(n2171), .B(n1598), .Z(mult_x_6_n1284) );
  AOI22_X1 U1793 ( .A1(mul_operand_b_q[23]), .A2(n628), .B1(
        mul_operand_b_q[22]), .B2(n606), .ZN(n1600) );
  AOI22_X1 U1794 ( .A1(mul_operand_b_q[21]), .A2(n2150), .B1(mult_x_6_n1081), 
        .B2(n1665), .ZN(n1599) );
  NAND2_X1 U1795 ( .A1(n1600), .A2(n1599), .ZN(n1601) );
  XOR2_X1 U1796 ( .A(n2171), .B(n1601), .Z(mult_x_6_n1285) );
  AOI22_X1 U1797 ( .A1(mul_operand_b_q[22]), .A2(n628), .B1(
        mul_operand_b_q[21]), .B2(n606), .ZN(n1603) );
  AOI22_X1 U1798 ( .A1(mul_operand_b_q[20]), .A2(n2150), .B1(mult_x_6_n1082), 
        .B2(n1665), .ZN(n1602) );
  NAND2_X1 U1799 ( .A1(n1603), .A2(n1602), .ZN(n1604) );
  XOR2_X1 U1800 ( .A(n2171), .B(n1604), .Z(mult_x_6_n1286) );
  AOI22_X1 U1801 ( .A1(mul_operand_b_q[21]), .A2(n628), .B1(
        mul_operand_b_q[20]), .B2(n606), .ZN(n1606) );
  AOI22_X1 U1802 ( .A1(mul_operand_b_q[19]), .A2(n2150), .B1(mult_x_6_n1083), 
        .B2(n1665), .ZN(n1605) );
  NAND2_X1 U1803 ( .A1(n1606), .A2(n1605), .ZN(n1607) );
  XOR2_X1 U1804 ( .A(n2171), .B(n1607), .Z(mult_x_6_n1287) );
  AOI22_X1 U1805 ( .A1(mul_operand_b_q[20]), .A2(n628), .B1(
        mul_operand_b_q[19]), .B2(n606), .ZN(n1609) );
  AOI22_X1 U1806 ( .A1(mul_operand_b_q[18]), .A2(n2150), .B1(mult_x_6_n1084), 
        .B2(n1665), .ZN(n1608) );
  NAND2_X1 U1807 ( .A1(n1609), .A2(n1608), .ZN(n1610) );
  XOR2_X1 U1808 ( .A(n2171), .B(n1610), .Z(mult_x_6_n1288) );
  AOI22_X1 U1809 ( .A1(mul_operand_b_q[19]), .A2(n628), .B1(
        mul_operand_b_q[18]), .B2(n606), .ZN(n1612) );
  AOI22_X1 U1810 ( .A1(mul_operand_b_q[17]), .A2(n2150), .B1(mult_x_6_n1085), 
        .B2(n1665), .ZN(n1611) );
  NAND2_X1 U1811 ( .A1(n1612), .A2(n1611), .ZN(n1613) );
  XOR2_X1 U1812 ( .A(n2171), .B(n1613), .Z(mult_x_6_n1289) );
  AOI22_X1 U1813 ( .A1(mul_operand_b_q[17]), .A2(n606), .B1(
        mul_operand_b_q[18]), .B2(n1666), .ZN(n1615) );
  AOI22_X1 U1814 ( .A1(n2185), .A2(n2150), .B1(mult_x_6_n1086), .B2(n1665), 
        .ZN(n1614) );
  NAND2_X1 U1815 ( .A1(n1615), .A2(n1614), .ZN(n1616) );
  XOR2_X1 U1816 ( .A(n2171), .B(n1616), .Z(mult_x_6_n1290) );
  AOI22_X1 U1817 ( .A1(mul_operand_b_q[17]), .A2(n628), .B1(n2184), .B2(n606), 
        .ZN(n1618) );
  AOI22_X1 U1818 ( .A1(mul_operand_b_q[15]), .A2(n2150), .B1(mult_x_6_n1087), 
        .B2(n1665), .ZN(n1617) );
  NAND2_X1 U1819 ( .A1(n1618), .A2(n1617), .ZN(n1619) );
  XOR2_X1 U1820 ( .A(n2171), .B(n1619), .Z(mult_x_6_n1291) );
  AOI22_X1 U1821 ( .A1(n2185), .A2(n628), .B1(mul_operand_b_q[15]), .B2(n606), 
        .ZN(n1621) );
  AOI22_X1 U1822 ( .A1(mul_operand_b_q[14]), .A2(n2150), .B1(mult_x_6_n1088), 
        .B2(n1665), .ZN(n1620) );
  NAND2_X1 U1823 ( .A1(n1621), .A2(n1620), .ZN(n1622) );
  XOR2_X1 U1824 ( .A(n2171), .B(n1622), .Z(mult_x_6_n1292) );
  AOI22_X1 U1825 ( .A1(mul_operand_b_q[15]), .A2(n628), .B1(
        mul_operand_b_q[14]), .B2(n606), .ZN(n1624) );
  AOI22_X1 U1826 ( .A1(mul_operand_b_q[13]), .A2(n2150), .B1(mult_x_6_n1089), 
        .B2(n1665), .ZN(n1623) );
  NAND2_X1 U1827 ( .A1(n1624), .A2(n1623), .ZN(n1625) );
  XOR2_X1 U1828 ( .A(n2171), .B(n1625), .Z(mult_x_6_n1293) );
  AOI22_X1 U1829 ( .A1(mul_operand_b_q[14]), .A2(n628), .B1(
        mul_operand_b_q[13]), .B2(n606), .ZN(n1627) );
  AOI22_X1 U1830 ( .A1(mul_operand_b_q[12]), .A2(n2150), .B1(mult_x_6_n1090), 
        .B2(n1665), .ZN(n1626) );
  NAND2_X1 U1831 ( .A1(n1627), .A2(n1626), .ZN(n1628) );
  XOR2_X1 U1832 ( .A(n2171), .B(n1628), .Z(mult_x_6_n1294) );
  AOI22_X1 U1833 ( .A1(mul_operand_b_q[13]), .A2(n628), .B1(
        mul_operand_b_q[12]), .B2(n606), .ZN(n1630) );
  AOI22_X1 U1834 ( .A1(mul_operand_b_q[11]), .A2(n2150), .B1(mult_x_6_n1091), 
        .B2(n1665), .ZN(n1629) );
  NAND2_X1 U1835 ( .A1(n1630), .A2(n1629), .ZN(n1631) );
  XOR2_X1 U1836 ( .A(n2171), .B(n1631), .Z(mult_x_6_n1295) );
  AOI22_X1 U1837 ( .A1(mul_operand_b_q[11]), .A2(n606), .B1(
        mul_operand_b_q[12]), .B2(n1666), .ZN(n1633) );
  AOI22_X1 U1838 ( .A1(mul_operand_b_q[10]), .A2(n2150), .B1(mult_x_6_n1092), 
        .B2(n1665), .ZN(n1632) );
  NAND2_X1 U1839 ( .A1(n1633), .A2(n1632), .ZN(n1634) );
  XOR2_X1 U1840 ( .A(n2171), .B(n1634), .Z(mult_x_6_n1296) );
  AOI22_X1 U1841 ( .A1(mul_operand_b_q[11]), .A2(n628), .B1(
        mul_operand_b_q[10]), .B2(n606), .ZN(n1636) );
  AOI22_X1 U1842 ( .A1(n2187), .A2(n2150), .B1(n2287), .B2(n1665), .ZN(n1635)
         );
  NAND2_X1 U1843 ( .A1(n1636), .A2(n1635), .ZN(n1637) );
  XOR2_X1 U1844 ( .A(n2171), .B(n1637), .Z(mult_x_6_n1297) );
  AOI22_X1 U1845 ( .A1(mul_operand_b_q[10]), .A2(n628), .B1(n2186), .B2(n606), 
        .ZN(n1639) );
  AOI22_X1 U1846 ( .A1(mul_operand_b_q[8]), .A2(n2150), .B1(mult_x_6_n1094), 
        .B2(n1665), .ZN(n1638) );
  NAND2_X1 U1847 ( .A1(n1639), .A2(n1638), .ZN(n1640) );
  XOR2_X1 U1848 ( .A(n2171), .B(n1640), .Z(mult_x_6_n1298) );
  AOI22_X1 U1849 ( .A1(n2187), .A2(n628), .B1(mul_operand_b_q[8]), .B2(n606), 
        .ZN(n1642) );
  AOI22_X1 U1850 ( .A1(mul_operand_b_q[7]), .A2(n2150), .B1(mult_x_6_n1095), 
        .B2(n1665), .ZN(n1641) );
  NAND2_X1 U1851 ( .A1(n1642), .A2(n1641), .ZN(n1643) );
  XOR2_X1 U1852 ( .A(n2171), .B(n1643), .Z(mult_x_6_n1299) );
  AOI22_X1 U1853 ( .A1(mul_operand_b_q[8]), .A2(n628), .B1(mul_operand_b_q[7]), 
        .B2(n606), .ZN(n1645) );
  AOI22_X1 U1854 ( .A1(n2189), .A2(n2150), .B1(mult_x_6_n1096), .B2(n1665), 
        .ZN(n1644) );
  NAND2_X1 U1855 ( .A1(n1645), .A2(n1644), .ZN(n1646) );
  XOR2_X1 U1856 ( .A(n2171), .B(n1646), .Z(mult_x_6_n1300) );
  AOI22_X1 U1857 ( .A1(mul_operand_b_q[7]), .A2(n628), .B1(n2188), .B2(n606), 
        .ZN(n1648) );
  AOI22_X1 U1858 ( .A1(n2191), .A2(n2150), .B1(n612), .B2(n1665), .ZN(n1647)
         );
  NAND2_X1 U1859 ( .A1(n1648), .A2(n1647), .ZN(n1649) );
  XOR2_X1 U1860 ( .A(n2171), .B(n1649), .Z(mult_x_6_n1301) );
  AOI22_X1 U1861 ( .A1(n2191), .A2(n606), .B1(n2188), .B2(n1666), .ZN(n1651)
         );
  AOI22_X1 U1862 ( .A1(mul_operand_b_q[4]), .A2(n2150), .B1(mult_x_6_n1098), 
        .B2(n1665), .ZN(n1650) );
  NAND2_X1 U1863 ( .A1(n1651), .A2(n1650), .ZN(n1652) );
  XOR2_X1 U1864 ( .A(n2171), .B(n1652), .Z(mult_x_6_n1302) );
  AOI22_X1 U1865 ( .A1(n2191), .A2(n628), .B1(n2192), .B2(n606), .ZN(n1654) );
  AOI22_X1 U1866 ( .A1(n2193), .A2(n2150), .B1(n355), .B2(n1665), .ZN(n1653)
         );
  NAND2_X1 U1867 ( .A1(n1654), .A2(n1653), .ZN(n1655) );
  XOR2_X1 U1868 ( .A(n2171), .B(n1655), .Z(mult_x_6_n1303) );
  AOI22_X1 U1869 ( .A1(mul_operand_b_q[4]), .A2(n628), .B1(n2193), .B2(n606), 
        .ZN(n1657) );
  AOI22_X1 U1870 ( .A1(n1009), .A2(n2150), .B1(n622), .B2(n1665), .ZN(n1656)
         );
  NAND2_X1 U1871 ( .A1(n1657), .A2(n1656), .ZN(n1658) );
  XOR2_X1 U1872 ( .A(n2171), .B(n1658), .Z(mult_x_6_n1304) );
  AOI22_X1 U1873 ( .A1(n2193), .A2(n628), .B1(n1009), .B2(n606), .ZN(n1660) );
  AOI22_X1 U1874 ( .A1(n2286), .A2(n2150), .B1(n833), .B2(n1665), .ZN(n1659)
         );
  NAND2_X1 U1875 ( .A1(n1660), .A2(n1659), .ZN(n1661) );
  XOR2_X1 U1876 ( .A(n2171), .B(n1661), .Z(mult_x_6_n1305) );
  AOI22_X1 U1877 ( .A1(n1009), .A2(n628), .B1(n2195), .B2(n606), .ZN(n1663) );
  AOI22_X1 U1878 ( .A1(n1018), .A2(n2150), .B1(mult_x_6_n1102), .B2(n1665), 
        .ZN(n1662) );
  NAND2_X1 U1879 ( .A1(n1663), .A2(n1662), .ZN(n1664) );
  XOR2_X1 U1880 ( .A(n2171), .B(n1664), .Z(mult_x_6_n1306) );
  XNOR2_X1 U1881 ( .A(mul_operand_a_q[11]), .B(mul_operand_a_q[12]), .ZN(n1670) );
  XOR2_X1 U1882 ( .A(mul_operand_a_q[14]), .B(mul_operand_a_q[13]), .Z(n1671)
         );
  XNOR2_X1 U1883 ( .A(mul_operand_a_q[13]), .B(mul_operand_a_q[12]), .ZN(n1667) );
  NAND3_X1 U1884 ( .A1(n1671), .A2(n1670), .A3(n1667), .ZN(n1672) );
  NAND3_X1 U1885 ( .A1(n1670), .A2(n1672), .A3(n2426), .ZN(n1668) );
  NAND2_X1 U1886 ( .A1(n1668), .A2(mul_operand_b_q[32]), .ZN(n1669) );
  XOR2_X1 U1887 ( .A(n2172), .B(n1669), .Z(mult_x_6_n1309) );
  NOR2_X1 U1888 ( .A1(n1670), .A2(n1671), .ZN(n1768) );
  OR2_X1 U1889 ( .A1(n2208), .A2(n2205), .ZN(n1673) );
  AOI222_X1 U1890 ( .A1(n1673), .A2(mul_operand_b_q[32]), .B1(mult_x_6_n1071), 
        .B2(n1767), .C1(n2179), .C2(n2148), .ZN(n1674) );
  XNOR2_X1 U1891 ( .A(n2172), .B(n1674), .ZN(mult_x_6_n1310) );
  AOI22_X1 U1892 ( .A1(n2180), .A2(n2148), .B1(mult_x_6_n1072), .B2(n1767), 
        .ZN(n1676) );
  NAND2_X1 U1893 ( .A1(n2177), .A2(n2208), .ZN(n1675) );
  OAI211_X1 U1894 ( .C1(n2178), .C2(n2426), .A(n1676), .B(n1675), .ZN(n1677)
         );
  XOR2_X1 U1895 ( .A(n2172), .B(n1677), .Z(mult_x_6_n1311) );
  AOI22_X1 U1896 ( .A1(n2179), .A2(n2208), .B1(n2180), .B2(n2205), .ZN(n1679)
         );
  AOI22_X1 U1897 ( .A1(mul_operand_b_q[29]), .A2(n2148), .B1(mult_x_6_n1073), 
        .B2(n1767), .ZN(n1678) );
  NAND2_X1 U1898 ( .A1(n1679), .A2(n1678), .ZN(n1680) );
  XOR2_X1 U1899 ( .A(n2172), .B(n1680), .Z(mult_x_6_n1312) );
  AOI22_X1 U1900 ( .A1(n2180), .A2(n2208), .B1(mul_operand_b_q[29]), .B2(n2205), .ZN(n1682) );
  AOI22_X1 U1901 ( .A1(n2181), .A2(n2148), .B1(mult_x_6_n1074), .B2(n1767), 
        .ZN(n1681) );
  NAND2_X1 U1902 ( .A1(n1682), .A2(n1681), .ZN(n1683) );
  XOR2_X1 U1903 ( .A(n2172), .B(n1683), .Z(mult_x_6_n1313) );
  AOI22_X1 U1904 ( .A1(mul_operand_b_q[29]), .A2(n2208), .B1(
        mul_operand_b_q[28]), .B2(n2205), .ZN(n1685) );
  AOI22_X1 U1905 ( .A1(mul_operand_b_q[27]), .A2(n2148), .B1(mult_x_6_n1075), 
        .B2(n1767), .ZN(n1684) );
  NAND2_X1 U1906 ( .A1(n1685), .A2(n1684), .ZN(n1686) );
  XOR2_X1 U1907 ( .A(n2172), .B(n1686), .Z(mult_x_6_n1314) );
  AOI22_X1 U1908 ( .A1(n2181), .A2(n6301), .B1(mul_operand_b_q[27]), .B2(n2205), .ZN(n1688) );
  AOI22_X1 U1909 ( .A1(n2182), .A2(n2148), .B1(mult_x_6_n1076), .B2(n1767), 
        .ZN(n1687) );
  NAND2_X1 U1910 ( .A1(n1688), .A2(n1687), .ZN(n1689) );
  XOR2_X1 U1911 ( .A(n2172), .B(n1689), .Z(mult_x_6_n1315) );
  AOI22_X1 U1912 ( .A1(mul_operand_b_q[27]), .A2(n6301), .B1(
        mul_operand_b_q[26]), .B2(n2205), .ZN(n1691) );
  AOI22_X1 U1913 ( .A1(mul_operand_b_q[25]), .A2(n2148), .B1(mult_x_6_n1077), 
        .B2(n1767), .ZN(n1690) );
  NAND2_X1 U1914 ( .A1(n1691), .A2(n1690), .ZN(n1692) );
  XOR2_X1 U1915 ( .A(n2172), .B(n1692), .Z(mult_x_6_n1316) );
  AOI22_X1 U1916 ( .A1(n2182), .A2(n6301), .B1(mul_operand_b_q[25]), .B2(n2205), .ZN(n1694) );
  AOI22_X1 U1917 ( .A1(n2183), .A2(n2148), .B1(mult_x_6_n1078), .B2(n1767), 
        .ZN(n1693) );
  NAND2_X1 U1918 ( .A1(n1694), .A2(n1693), .ZN(n1695) );
  XOR2_X1 U1919 ( .A(n2172), .B(n1695), .Z(mult_x_6_n1317) );
  AOI22_X1 U1920 ( .A1(mul_operand_b_q[25]), .A2(n6301), .B1(
        mul_operand_b_q[24]), .B2(n2206), .ZN(n1697) );
  AOI22_X1 U1921 ( .A1(mul_operand_b_q[23]), .A2(n2148), .B1(mult_x_6_n1079), 
        .B2(n1767), .ZN(n1696) );
  NAND2_X1 U1922 ( .A1(n1697), .A2(n1696), .ZN(n1698) );
  XOR2_X1 U1923 ( .A(n2172), .B(n1698), .Z(mult_x_6_n1318) );
  AOI22_X1 U1924 ( .A1(n2183), .A2(n6301), .B1(mul_operand_b_q[23]), .B2(n2206), .ZN(n17001) );
  AOI22_X1 U1925 ( .A1(mul_operand_b_q[22]), .A2(n2148), .B1(mult_x_6_n1080), 
        .B2(n1767), .ZN(n1699) );
  NAND2_X1 U1926 ( .A1(n17001), .A2(n1699), .ZN(n1701) );
  XOR2_X1 U1927 ( .A(n2172), .B(n1701), .Z(mult_x_6_n1319) );
  AOI22_X1 U1928 ( .A1(mul_operand_b_q[23]), .A2(n6301), .B1(
        mul_operand_b_q[22]), .B2(n2206), .ZN(n1703) );
  AOI22_X1 U1929 ( .A1(mul_operand_b_q[21]), .A2(n2148), .B1(mult_x_6_n1081), 
        .B2(n1767), .ZN(n1702) );
  NAND2_X1 U1930 ( .A1(n1703), .A2(n1702), .ZN(n1704) );
  XOR2_X1 U1931 ( .A(n2172), .B(n1704), .Z(mult_x_6_n1320) );
  AOI22_X1 U1932 ( .A1(mul_operand_b_q[22]), .A2(n6301), .B1(
        mul_operand_b_q[21]), .B2(n2206), .ZN(n1706) );
  AOI22_X1 U1933 ( .A1(mul_operand_b_q[20]), .A2(n2148), .B1(mult_x_6_n1082), 
        .B2(n1767), .ZN(n1705) );
  NAND2_X1 U1934 ( .A1(n1706), .A2(n1705), .ZN(n1707) );
  XOR2_X1 U1935 ( .A(n2172), .B(n1707), .Z(mult_x_6_n1321) );
  AOI22_X1 U1936 ( .A1(mul_operand_b_q[21]), .A2(n6301), .B1(
        mul_operand_b_q[20]), .B2(n2206), .ZN(n1709) );
  AOI22_X1 U1937 ( .A1(mul_operand_b_q[19]), .A2(n2148), .B1(mult_x_6_n1083), 
        .B2(n1767), .ZN(n1708) );
  NAND2_X1 U1938 ( .A1(n1709), .A2(n1708), .ZN(n17101) );
  XOR2_X1 U1939 ( .A(n2172), .B(n17101), .Z(mult_x_6_n1322) );
  AOI22_X1 U1940 ( .A1(mul_operand_b_q[20]), .A2(n6301), .B1(
        mul_operand_b_q[19]), .B2(n2206), .ZN(n1712) );
  AOI22_X1 U1941 ( .A1(mul_operand_b_q[18]), .A2(n2148), .B1(mult_x_6_n1084), 
        .B2(n1767), .ZN(n1711) );
  NAND2_X1 U1942 ( .A1(n1712), .A2(n1711), .ZN(n1713) );
  XOR2_X1 U1943 ( .A(n2172), .B(n1713), .Z(mult_x_6_n1323) );
  AOI22_X1 U1944 ( .A1(mul_operand_b_q[19]), .A2(n6301), .B1(
        mul_operand_b_q[18]), .B2(n2206), .ZN(n1715) );
  AOI22_X1 U1945 ( .A1(mul_operand_b_q[17]), .A2(n2148), .B1(mult_x_6_n1085), 
        .B2(n1767), .ZN(n1714) );
  NAND2_X1 U1946 ( .A1(n1715), .A2(n1714), .ZN(n1716) );
  XOR2_X1 U1947 ( .A(n2172), .B(n1716), .Z(mult_x_6_n1324) );
  AOI22_X1 U1948 ( .A1(mul_operand_b_q[17]), .A2(n2207), .B1(
        mul_operand_b_q[18]), .B2(n2208), .ZN(n1718) );
  AOI22_X1 U1949 ( .A1(n2185), .A2(n2148), .B1(mult_x_6_n1086), .B2(n1767), 
        .ZN(n1717) );
  NAND2_X1 U1950 ( .A1(n1718), .A2(n1717), .ZN(n1719) );
  XOR2_X1 U1951 ( .A(n2172), .B(n1719), .Z(mult_x_6_n1325) );
  AOI22_X1 U1952 ( .A1(mul_operand_b_q[17]), .A2(n6301), .B1(n2184), .B2(n2206), .ZN(n1721) );
  AOI22_X1 U1953 ( .A1(mul_operand_b_q[15]), .A2(n2148), .B1(mult_x_6_n1087), 
        .B2(n1767), .ZN(n17201) );
  NAND2_X1 U1954 ( .A1(n1721), .A2(n17201), .ZN(n1722) );
  XOR2_X1 U1955 ( .A(n2172), .B(n1722), .Z(mult_x_6_n1326) );
  AOI22_X1 U1956 ( .A1(n2185), .A2(n6301), .B1(mul_operand_b_q[15]), .B2(n2206), .ZN(n1724) );
  AOI22_X1 U1957 ( .A1(mul_operand_b_q[14]), .A2(n2148), .B1(mult_x_6_n1088), 
        .B2(n1767), .ZN(n1723) );
  NAND2_X1 U1958 ( .A1(n1724), .A2(n1723), .ZN(n1725) );
  XOR2_X1 U1959 ( .A(n2172), .B(n1725), .Z(mult_x_6_n1327) );
  AOI22_X1 U1960 ( .A1(mul_operand_b_q[15]), .A2(n6301), .B1(
        mul_operand_b_q[14]), .B2(n2206), .ZN(n1727) );
  AOI22_X1 U1961 ( .A1(mul_operand_b_q[13]), .A2(n2148), .B1(mult_x_6_n1089), 
        .B2(n1767), .ZN(n1726) );
  NAND2_X1 U1962 ( .A1(n1727), .A2(n1726), .ZN(n1728) );
  XOR2_X1 U1963 ( .A(n2172), .B(n1728), .Z(mult_x_6_n1328) );
  AOI22_X1 U1964 ( .A1(mul_operand_b_q[14]), .A2(n6301), .B1(
        mul_operand_b_q[13]), .B2(n2207), .ZN(n17301) );
  AOI22_X1 U1965 ( .A1(mul_operand_b_q[12]), .A2(n2148), .B1(mult_x_6_n1090), 
        .B2(n2204), .ZN(n1729) );
  NAND2_X1 U1966 ( .A1(n17301), .A2(n1729), .ZN(n1731) );
  XOR2_X1 U1967 ( .A(n2172), .B(n1731), .Z(mult_x_6_n1329) );
  AOI22_X1 U1968 ( .A1(mul_operand_b_q[13]), .A2(n6301), .B1(
        mul_operand_b_q[12]), .B2(n2207), .ZN(n1733) );
  AOI22_X1 U1969 ( .A1(mul_operand_b_q[11]), .A2(n2148), .B1(mult_x_6_n1091), 
        .B2(n2204), .ZN(n1732) );
  NAND2_X1 U1970 ( .A1(n1733), .A2(n1732), .ZN(n1734) );
  XOR2_X1 U1971 ( .A(n2172), .B(n1734), .Z(mult_x_6_n1330) );
  AOI22_X1 U1972 ( .A1(mul_operand_b_q[11]), .A2(n2207), .B1(
        mul_operand_b_q[12]), .B2(n2208), .ZN(n1736) );
  AOI22_X1 U1973 ( .A1(mul_operand_b_q[10]), .A2(n2148), .B1(mult_x_6_n1092), 
        .B2(n2204), .ZN(n1735) );
  NAND2_X1 U1974 ( .A1(n1736), .A2(n1735), .ZN(n1737) );
  XOR2_X1 U1975 ( .A(n2172), .B(n1737), .Z(mult_x_6_n1331) );
  AOI22_X1 U1976 ( .A1(mul_operand_b_q[11]), .A2(n6301), .B1(
        mul_operand_b_q[10]), .B2(n2206), .ZN(n1739) );
  AOI22_X1 U1977 ( .A1(n2187), .A2(n2148), .B1(n2287), .B2(n2204), .ZN(n1738)
         );
  NAND2_X1 U1978 ( .A1(n1739), .A2(n1738), .ZN(n17401) );
  XOR2_X1 U1979 ( .A(n2172), .B(n17401), .Z(mult_x_6_n1332) );
  AOI22_X1 U1980 ( .A1(mul_operand_b_q[10]), .A2(n6301), .B1(n2186), .B2(n2207), .ZN(n1742) );
  AOI22_X1 U1981 ( .A1(mul_operand_b_q[8]), .A2(n2148), .B1(mult_x_6_n1094), 
        .B2(n2204), .ZN(n1741) );
  NAND2_X1 U1982 ( .A1(n1742), .A2(n1741), .ZN(n1743) );
  XOR2_X1 U1983 ( .A(n2172), .B(n1743), .Z(mult_x_6_n1333) );
  AOI22_X1 U1984 ( .A1(n2187), .A2(n6301), .B1(mul_operand_b_q[8]), .B2(n2206), 
        .ZN(n1745) );
  AOI22_X1 U1985 ( .A1(mul_operand_b_q[7]), .A2(n2148), .B1(mult_x_6_n1095), 
        .B2(n2204), .ZN(n1744) );
  NAND2_X1 U1986 ( .A1(n1745), .A2(n1744), .ZN(n1746) );
  XOR2_X1 U1987 ( .A(n2172), .B(n1746), .Z(mult_x_6_n1334) );
  AOI22_X1 U1988 ( .A1(mul_operand_b_q[8]), .A2(n6301), .B1(mul_operand_b_q[7]), .B2(n2207), .ZN(n1748) );
  AOI22_X1 U1989 ( .A1(n2189), .A2(n2148), .B1(mult_x_6_n1096), .B2(n2204), 
        .ZN(n1747) );
  NAND2_X1 U1990 ( .A1(n1748), .A2(n1747), .ZN(n1749) );
  XOR2_X1 U1991 ( .A(n2172), .B(n1749), .Z(mult_x_6_n1335) );
  AOI22_X1 U1992 ( .A1(mul_operand_b_q[7]), .A2(n6301), .B1(n2188), .B2(n2207), 
        .ZN(n1751) );
  AOI22_X1 U1993 ( .A1(n2191), .A2(n2148), .B1(n612), .B2(n2204), .ZN(n17501)
         );
  NAND2_X1 U1994 ( .A1(n1751), .A2(n17501), .ZN(n1752) );
  XOR2_X1 U1995 ( .A(n2172), .B(n1752), .Z(mult_x_6_n1336) );
  AOI22_X1 U1996 ( .A1(n2191), .A2(n2207), .B1(n2188), .B2(n2208), .ZN(n1754)
         );
  AOI22_X1 U1997 ( .A1(mul_operand_b_q[4]), .A2(n2148), .B1(mult_x_6_n1098), 
        .B2(n2204), .ZN(n1753) );
  NAND2_X1 U1998 ( .A1(n1754), .A2(n1753), .ZN(n1755) );
  XOR2_X1 U1999 ( .A(n2172), .B(n1755), .Z(mult_x_6_n1337) );
  AOI22_X1 U2000 ( .A1(n2191), .A2(n6301), .B1(n2192), .B2(n2207), .ZN(n1757)
         );
  AOI22_X1 U2001 ( .A1(n2193), .A2(n2148), .B1(n355), .B2(n2204), .ZN(n1756)
         );
  NAND2_X1 U2002 ( .A1(n1757), .A2(n1756), .ZN(n1758) );
  XOR2_X1 U2003 ( .A(n2172), .B(n1758), .Z(mult_x_6_n1338) );
  AOI22_X1 U2004 ( .A1(mul_operand_b_q[4]), .A2(n6301), .B1(n2193), .B2(n2207), 
        .ZN(n17601) );
  AOI22_X1 U2005 ( .A1(n1009), .A2(n2148), .B1(n622), .B2(n2204), .ZN(n1759)
         );
  NAND2_X1 U2006 ( .A1(n17601), .A2(n1759), .ZN(n1761) );
  XOR2_X1 U2007 ( .A(n2172), .B(n1761), .Z(mult_x_6_n1339) );
  AOI22_X1 U2008 ( .A1(n2193), .A2(n6301), .B1(n1009), .B2(n2207), .ZN(n1762)
         );
  XOR2_X1 U2009 ( .A(n2172), .B(n1763), .Z(mult_x_6_n1340) );
  AOI22_X1 U2010 ( .A1(n1009), .A2(n6301), .B1(n2286), .B2(n2207), .ZN(n1765)
         );
  AOI22_X1 U2011 ( .A1(n2196), .A2(n2148), .B1(mult_x_6_n1102), .B2(n2204), 
        .ZN(n1764) );
  NAND2_X1 U2012 ( .A1(n1765), .A2(n1764), .ZN(n1766) );
  XOR2_X1 U2013 ( .A(n2172), .B(n1766), .Z(mult_x_6_n1341) );
  XNOR2_X1 U2014 ( .A(mul_operand_a_q[8]), .B(mul_operand_a_q[9]), .ZN(n1772)
         );
  XOR2_X1 U2015 ( .A(mul_operand_a_q[11]), .B(mul_operand_a_q[10]), .Z(n1773)
         );
  XNOR2_X1 U2016 ( .A(mul_operand_a_q[10]), .B(mul_operand_a_q[9]), .ZN(n1769)
         );
  NAND3_X1 U2017 ( .A1(n1773), .A2(n1772), .A3(n1769), .ZN(n1774) );
  NAND3_X1 U2018 ( .A1(n1772), .A2(n1774), .A3(n2210), .ZN(n17701) );
  NAND2_X1 U2019 ( .A1(n17701), .A2(mul_operand_b_q[32]), .ZN(n1771) );
  XOR2_X1 U2020 ( .A(n2173), .B(n1771), .Z(mult_x_6_n1344) );
  NOR2_X1 U2021 ( .A1(n1772), .A2(n1773), .ZN(n1869) );
  OR2_X1 U2022 ( .A1(n2212), .A2(n2211), .ZN(n1775) );
  AOI222_X1 U2023 ( .A1(n1775), .A2(mul_operand_b_q[32]), .B1(mult_x_6_n1071), 
        .B2(n1868), .C1(n2179), .C2(n2146), .ZN(n1776) );
  XNOR2_X1 U2024 ( .A(n2173), .B(n1776), .ZN(mult_x_6_n1345) );
  AOI22_X1 U2025 ( .A1(n2180), .A2(n2146), .B1(mult_x_6_n1072), .B2(n1868), 
        .ZN(n1778) );
  NAND2_X1 U2026 ( .A1(n2177), .A2(n2212), .ZN(n1777) );
  OAI211_X1 U2027 ( .C1(n2178), .C2(n2210), .A(n1778), .B(n1777), .ZN(n1779)
         );
  XOR2_X1 U2028 ( .A(n2173), .B(n1779), .Z(mult_x_6_n1346) );
  AOI22_X1 U2029 ( .A1(n2180), .A2(n2211), .B1(mul_operand_b_q[29]), .B2(n2146), .ZN(n1781) );
  AOI22_X1 U2030 ( .A1(n2179), .A2(n2212), .B1(mult_x_6_n1073), .B2(n1868), 
        .ZN(n17801) );
  NAND2_X1 U2031 ( .A1(n1781), .A2(n17801), .ZN(n1782) );
  XOR2_X1 U2032 ( .A(n2173), .B(n1782), .Z(mult_x_6_n1347) );
  AOI22_X1 U2033 ( .A1(n2180), .A2(n2212), .B1(mul_operand_b_q[28]), .B2(n2146), .ZN(n1784) );
  AOI22_X1 U2034 ( .A1(mul_operand_b_q[29]), .A2(n2211), .B1(mult_x_6_n1074), 
        .B2(n1868), .ZN(n1783) );
  NAND2_X1 U2035 ( .A1(n1784), .A2(n1783), .ZN(n1785) );
  XOR2_X1 U2036 ( .A(n2173), .B(n1785), .Z(mult_x_6_n1348) );
  AOI22_X1 U2037 ( .A1(mul_operand_b_q[29]), .A2(n2212), .B1(
        mul_operand_b_q[27]), .B2(n2146), .ZN(n1787) );
  AOI22_X1 U2038 ( .A1(n2181), .A2(n2211), .B1(mult_x_6_n1075), .B2(n1868), 
        .ZN(n1786) );
  NAND2_X1 U2039 ( .A1(n1787), .A2(n1786), .ZN(n1788) );
  XOR2_X1 U2040 ( .A(n2173), .B(n1788), .Z(mult_x_6_n1349) );
  AOI22_X1 U2041 ( .A1(n2181), .A2(n2212), .B1(mul_operand_b_q[26]), .B2(n2146), .ZN(n17901) );
  AOI22_X1 U2042 ( .A1(mul_operand_b_q[27]), .A2(n2211), .B1(mult_x_6_n1076), 
        .B2(n1868), .ZN(n1789) );
  NAND2_X1 U2043 ( .A1(n17901), .A2(n1789), .ZN(n1791) );
  XOR2_X1 U2044 ( .A(n2173), .B(n1791), .Z(mult_x_6_n1350) );
  AOI22_X1 U2045 ( .A1(mul_operand_b_q[27]), .A2(n2212), .B1(
        mul_operand_b_q[25]), .B2(n2146), .ZN(n1793) );
  AOI22_X1 U2046 ( .A1(n2182), .A2(n2211), .B1(mult_x_6_n1077), .B2(n1868), 
        .ZN(n1792) );
  NAND2_X1 U2047 ( .A1(n1793), .A2(n1792), .ZN(n1794) );
  XOR2_X1 U2048 ( .A(n2173), .B(n1794), .Z(mult_x_6_n1351) );
  AOI22_X1 U2049 ( .A1(n2182), .A2(n2212), .B1(mul_operand_b_q[24]), .B2(n2146), .ZN(n1796) );
  AOI22_X1 U2050 ( .A1(mul_operand_b_q[25]), .A2(n2211), .B1(mult_x_6_n1078), 
        .B2(n1868), .ZN(n1795) );
  NAND2_X1 U2051 ( .A1(n1796), .A2(n1795), .ZN(n1797) );
  XOR2_X1 U2052 ( .A(n2173), .B(n1797), .Z(mult_x_6_n1352) );
  AOI22_X1 U2053 ( .A1(mul_operand_b_q[25]), .A2(n629), .B1(
        mul_operand_b_q[23]), .B2(n2146), .ZN(n1799) );
  AOI22_X1 U2054 ( .A1(n2183), .A2(n602), .B1(mult_x_6_n1079), .B2(n2209), 
        .ZN(n1798) );
  NAND2_X1 U2055 ( .A1(n1799), .A2(n1798), .ZN(n18001) );
  XOR2_X1 U2056 ( .A(n2173), .B(n18001), .Z(mult_x_6_n1353) );
  AOI22_X1 U2057 ( .A1(n2183), .A2(n629), .B1(mul_operand_b_q[22]), .B2(n2146), 
        .ZN(n1802) );
  AOI22_X1 U2058 ( .A1(mul_operand_b_q[23]), .A2(n602), .B1(mult_x_6_n1080), 
        .B2(n2209), .ZN(n1801) );
  NAND2_X1 U2059 ( .A1(n1802), .A2(n1801), .ZN(n1803) );
  XOR2_X1 U2060 ( .A(n2173), .B(n1803), .Z(mult_x_6_n1354) );
  AOI22_X1 U2061 ( .A1(mul_operand_b_q[23]), .A2(n629), .B1(
        mul_operand_b_q[21]), .B2(n2146), .ZN(n1805) );
  AOI22_X1 U2062 ( .A1(mul_operand_b_q[22]), .A2(n602), .B1(mult_x_6_n1081), 
        .B2(n2209), .ZN(n1804) );
  NAND2_X1 U2063 ( .A1(n1805), .A2(n1804), .ZN(n1806) );
  XOR2_X1 U2064 ( .A(n2173), .B(n1806), .Z(mult_x_6_n1355) );
  AOI22_X1 U2065 ( .A1(mul_operand_b_q[22]), .A2(n629), .B1(
        mul_operand_b_q[20]), .B2(n2146), .ZN(n1808) );
  AOI22_X1 U2066 ( .A1(mul_operand_b_q[21]), .A2(n602), .B1(mult_x_6_n1082), 
        .B2(n2209), .ZN(n1807) );
  NAND2_X1 U2067 ( .A1(n1808), .A2(n1807), .ZN(n1809) );
  XOR2_X1 U2068 ( .A(n2173), .B(n1809), .Z(mult_x_6_n1356) );
  AOI22_X1 U2069 ( .A1(mul_operand_b_q[21]), .A2(n629), .B1(
        mul_operand_b_q[19]), .B2(n2146), .ZN(n1811) );
  AOI22_X1 U2070 ( .A1(mul_operand_b_q[20]), .A2(n602), .B1(mult_x_6_n1083), 
        .B2(n2209), .ZN(n18101) );
  NAND2_X1 U2071 ( .A1(n1811), .A2(n18101), .ZN(n1812) );
  XOR2_X1 U2072 ( .A(n2173), .B(n1812), .Z(mult_x_6_n1357) );
  AOI22_X1 U2073 ( .A1(mul_operand_b_q[20]), .A2(n629), .B1(
        mul_operand_b_q[18]), .B2(n2146), .ZN(n1814) );
  AOI22_X1 U2074 ( .A1(mul_operand_b_q[19]), .A2(n602), .B1(mult_x_6_n1084), 
        .B2(n2209), .ZN(n1813) );
  NAND2_X1 U2075 ( .A1(n1814), .A2(n1813), .ZN(n1815) );
  XOR2_X1 U2076 ( .A(n2173), .B(n1815), .Z(mult_x_6_n1358) );
  AOI22_X1 U2077 ( .A1(mul_operand_b_q[19]), .A2(n629), .B1(
        mul_operand_b_q[17]), .B2(n2146), .ZN(n1817) );
  AOI22_X1 U2078 ( .A1(mul_operand_b_q[18]), .A2(n602), .B1(mult_x_6_n1085), 
        .B2(n2209), .ZN(n1816) );
  NAND2_X1 U2079 ( .A1(n1817), .A2(n1816), .ZN(n1818) );
  XOR2_X1 U2080 ( .A(n2173), .B(n1818), .Z(mult_x_6_n1359) );
  AOI22_X1 U2081 ( .A1(mul_operand_b_q[18]), .A2(n629), .B1(n2184), .B2(n2146), 
        .ZN(n18201) );
  AOI22_X1 U2082 ( .A1(mul_operand_b_q[17]), .A2(n602), .B1(mult_x_6_n1086), 
        .B2(n2209), .ZN(n1819) );
  NAND2_X1 U2083 ( .A1(n18201), .A2(n1819), .ZN(n1821) );
  XOR2_X1 U2084 ( .A(n2173), .B(n1821), .Z(mult_x_6_n1360) );
  AOI22_X1 U2085 ( .A1(mul_operand_b_q[17]), .A2(n629), .B1(
        mul_operand_b_q[15]), .B2(n2146), .ZN(n1823) );
  AOI22_X1 U2086 ( .A1(n2185), .A2(n602), .B1(mult_x_6_n1087), .B2(n2209), 
        .ZN(n1822) );
  NAND2_X1 U2087 ( .A1(n1823), .A2(n1822), .ZN(n1824) );
  XOR2_X1 U2088 ( .A(n2173), .B(n1824), .Z(mult_x_6_n1361) );
  AOI22_X1 U2089 ( .A1(n2185), .A2(n629), .B1(mul_operand_b_q[14]), .B2(n2146), 
        .ZN(n1826) );
  AOI22_X1 U2090 ( .A1(mul_operand_b_q[15]), .A2(n602), .B1(mult_x_6_n1088), 
        .B2(n2209), .ZN(n1825) );
  NAND2_X1 U2091 ( .A1(n1826), .A2(n1825), .ZN(n1827) );
  XOR2_X1 U2092 ( .A(n2173), .B(n1827), .Z(mult_x_6_n1362) );
  AOI22_X1 U2093 ( .A1(mul_operand_b_q[15]), .A2(n629), .B1(
        mul_operand_b_q[13]), .B2(n2146), .ZN(n1829) );
  AOI22_X1 U2094 ( .A1(mul_operand_b_q[14]), .A2(n602), .B1(mult_x_6_n1089), 
        .B2(n2209), .ZN(n1828) );
  NAND2_X1 U2095 ( .A1(n1829), .A2(n1828), .ZN(n18301) );
  XOR2_X1 U2096 ( .A(n2173), .B(n18301), .Z(mult_x_6_n1363) );
  AOI22_X1 U2097 ( .A1(mul_operand_b_q[14]), .A2(n629), .B1(
        mul_operand_b_q[12]), .B2(n2146), .ZN(n1832) );
  AOI22_X1 U2098 ( .A1(mul_operand_b_q[13]), .A2(n602), .B1(mult_x_6_n1090), 
        .B2(n1868), .ZN(n1831) );
  NAND2_X1 U2099 ( .A1(n1832), .A2(n1831), .ZN(n1833) );
  XOR2_X1 U2100 ( .A(n2173), .B(n1833), .Z(mult_x_6_n1364) );
  AOI22_X1 U2101 ( .A1(mul_operand_b_q[13]), .A2(n629), .B1(
        mul_operand_b_q[11]), .B2(n2146), .ZN(n1835) );
  AOI22_X1 U2102 ( .A1(mul_operand_b_q[12]), .A2(n602), .B1(mult_x_6_n1091), 
        .B2(n1868), .ZN(n1834) );
  NAND2_X1 U2103 ( .A1(n1835), .A2(n1834), .ZN(n1836) );
  XOR2_X1 U2104 ( .A(n2173), .B(n1836), .Z(mult_x_6_n1365) );
  AOI22_X1 U2105 ( .A1(mul_operand_b_q[12]), .A2(n629), .B1(
        mul_operand_b_q[10]), .B2(n2146), .ZN(n1838) );
  AOI22_X1 U2106 ( .A1(mul_operand_b_q[11]), .A2(n602), .B1(mult_x_6_n1092), 
        .B2(n1868), .ZN(n1837) );
  NAND2_X1 U2107 ( .A1(n1838), .A2(n1837), .ZN(n1839) );
  XOR2_X1 U2108 ( .A(n2173), .B(n1839), .Z(mult_x_6_n1366) );
  AOI22_X1 U2109 ( .A1(mul_operand_b_q[11]), .A2(n629), .B1(n2186), .B2(n2146), 
        .ZN(n1841) );
  AOI22_X1 U2110 ( .A1(mul_operand_b_q[10]), .A2(n602), .B1(n2287), .B2(n1868), 
        .ZN(n18401) );
  NAND2_X1 U2111 ( .A1(n1841), .A2(n18401), .ZN(n1842) );
  XOR2_X1 U2112 ( .A(n2173), .B(n1842), .Z(mult_x_6_n1367) );
  AOI22_X1 U2113 ( .A1(mul_operand_b_q[10]), .A2(n629), .B1(mul_operand_b_q[8]), .B2(n2146), .ZN(n1844) );
  AOI22_X1 U2114 ( .A1(n2187), .A2(n602), .B1(mult_x_6_n1094), .B2(n1868), 
        .ZN(n1843) );
  NAND2_X1 U2115 ( .A1(n1844), .A2(n1843), .ZN(n1845) );
  XOR2_X1 U2116 ( .A(n2173), .B(n1845), .Z(mult_x_6_n1368) );
  AOI22_X1 U2117 ( .A1(n2187), .A2(n629), .B1(mul_operand_b_q[7]), .B2(n2146), 
        .ZN(n1847) );
  AOI22_X1 U2118 ( .A1(mul_operand_b_q[8]), .A2(n602), .B1(mult_x_6_n1095), 
        .B2(n2209), .ZN(n1846) );
  NAND2_X1 U2119 ( .A1(n1847), .A2(n1846), .ZN(n1848) );
  XOR2_X1 U2120 ( .A(n2173), .B(n1848), .Z(mult_x_6_n1369) );
  AOI22_X1 U2121 ( .A1(mul_operand_b_q[8]), .A2(n629), .B1(n2188), .B2(n2146), 
        .ZN(n18501) );
  AOI22_X1 U2122 ( .A1(mul_operand_b_q[7]), .A2(n602), .B1(mult_x_6_n1096), 
        .B2(n2209), .ZN(n1849) );
  NAND2_X1 U2123 ( .A1(n18501), .A2(n1849), .ZN(n1851) );
  XOR2_X1 U2124 ( .A(n2173), .B(n1851), .Z(mult_x_6_n1370) );
  AOI22_X1 U2125 ( .A1(mul_operand_b_q[7]), .A2(n629), .B1(n2190), .B2(n2146), 
        .ZN(n1853) );
  AOI22_X1 U2126 ( .A1(n2189), .A2(n602), .B1(n612), .B2(n1868), .ZN(n1852) );
  NAND2_X1 U2127 ( .A1(n1853), .A2(n1852), .ZN(n1854) );
  XOR2_X1 U2128 ( .A(n2173), .B(n1854), .Z(mult_x_6_n1371) );
  AOI22_X1 U2129 ( .A1(n2189), .A2(n629), .B1(n2192), .B2(n2146), .ZN(n1856)
         );
  AOI22_X1 U2130 ( .A1(n2190), .A2(n602), .B1(mult_x_6_n1098), .B2(n1868), 
        .ZN(n1855) );
  NAND2_X1 U2131 ( .A1(n1856), .A2(n1855), .ZN(n1857) );
  XOR2_X1 U2132 ( .A(n2173), .B(n1857), .Z(mult_x_6_n1372) );
  AOI22_X1 U2133 ( .A1(n2190), .A2(n629), .B1(n2193), .B2(n2146), .ZN(n1859)
         );
  AOI22_X1 U2134 ( .A1(mul_operand_b_q[4]), .A2(n602), .B1(n355), .B2(n2209), 
        .ZN(n1858) );
  NAND2_X1 U2135 ( .A1(n1859), .A2(n1858), .ZN(n18601) );
  XOR2_X1 U2136 ( .A(n2173), .B(n18601), .Z(mult_x_6_n1373) );
  AOI22_X1 U2137 ( .A1(mul_operand_b_q[4]), .A2(n629), .B1(n1009), .B2(n2146), 
        .ZN(n1862) );
  AOI22_X1 U2138 ( .A1(n2193), .A2(n602), .B1(n622), .B2(n2209), .ZN(n1861) );
  AOI22_X1 U2139 ( .A1(n2193), .A2(n629), .B1(n2195), .B2(n2146), .ZN(n1863)
         );
  XOR2_X1 U2140 ( .A(n2173), .B(n1864), .Z(mult_x_6_n1375) );
  AOI22_X1 U2141 ( .A1(n1009), .A2(n629), .B1(n2196), .B2(n2146), .ZN(n1866)
         );
  AOI22_X1 U2142 ( .A1(n2286), .A2(n602), .B1(mult_x_6_n1102), .B2(n2209), 
        .ZN(n1865) );
  NAND2_X1 U2143 ( .A1(n1866), .A2(n1865), .ZN(n1867) );
  XOR2_X1 U2144 ( .A(n2173), .B(n1867), .Z(mult_x_6_n1376) );
  XNOR2_X1 U2145 ( .A(mul_operand_a_q[7]), .B(mul_operand_a_q[6]), .ZN(n18701)
         );
  NAND3_X1 U2146 ( .A1(n1874), .A2(n18701), .A3(n1873), .ZN(n1875) );
  NAND3_X1 U2147 ( .A1(n1873), .A2(n1875), .A3(n2215), .ZN(n1871) );
  NAND2_X1 U2148 ( .A1(n1871), .A2(n2177), .ZN(n1872) );
  XOR2_X1 U2149 ( .A(n2174), .B(n1872), .Z(mult_x_6_n1379) );
  OR2_X1 U2150 ( .A1(n2218), .A2(n1020), .ZN(n1876) );
  AOI222_X1 U2151 ( .A1(n1876), .A2(mul_operand_b_q[32]), .B1(mult_x_6_n1071), 
        .B2(n2213), .C1(n2179), .C2(n2226), .ZN(n1877) );
  XNOR2_X1 U2152 ( .A(n2174), .B(n1877), .ZN(mult_x_6_n1380) );
  AOI22_X1 U2153 ( .A1(n2180), .A2(n405), .B1(mult_x_6_n1072), .B2(n2213), 
        .ZN(n1879) );
  NAND2_X1 U2154 ( .A1(n2177), .A2(n2217), .ZN(n1878) );
  OAI211_X1 U2155 ( .C1(n2178), .C2(n2215), .A(n1879), .B(n1878), .ZN(n18801)
         );
  XOR2_X1 U2156 ( .A(n2174), .B(n18801), .Z(mult_x_6_n1381) );
  AOI22_X1 U2157 ( .A1(n2179), .A2(n2218), .B1(n2180), .B2(n1020), .ZN(n1882)
         );
  AOI22_X1 U2158 ( .A1(mul_operand_b_q[29]), .A2(n405), .B1(mult_x_6_n1073), 
        .B2(n2213), .ZN(n1881) );
  NAND2_X1 U2159 ( .A1(n1882), .A2(n1881), .ZN(n1883) );
  XOR2_X1 U2160 ( .A(n2174), .B(n1883), .Z(mult_x_6_n1382) );
  AOI22_X1 U2161 ( .A1(n2180), .A2(n2217), .B1(mul_operand_b_q[29]), .B2(n1020), .ZN(n1885) );
  AOI22_X1 U2162 ( .A1(n2181), .A2(n2226), .B1(mult_x_6_n1074), .B2(n2213), 
        .ZN(n1884) );
  NAND2_X1 U2163 ( .A1(n1885), .A2(n1884), .ZN(n1886) );
  XOR2_X1 U2164 ( .A(n2174), .B(n1886), .Z(mult_x_6_n1383) );
  AOI22_X1 U2165 ( .A1(mul_operand_b_q[29]), .A2(n2218), .B1(
        mul_operand_b_q[28]), .B2(n1020), .ZN(n1888) );
  AOI22_X1 U2166 ( .A1(mul_operand_b_q[27]), .A2(n405), .B1(mult_x_6_n1075), 
        .B2(n2213), .ZN(n1887) );
  NAND2_X1 U2167 ( .A1(n1888), .A2(n1887), .ZN(n1889) );
  XOR2_X1 U2168 ( .A(n2174), .B(n1889), .Z(mult_x_6_n1384) );
  AOI22_X1 U2169 ( .A1(n2181), .A2(n2217), .B1(mul_operand_b_q[27]), .B2(n1020), .ZN(n1891) );
  AOI22_X1 U2170 ( .A1(n2182), .A2(n405), .B1(mult_x_6_n1076), .B2(n2213), 
        .ZN(n18901) );
  NAND2_X1 U2171 ( .A1(n1891), .A2(n18901), .ZN(n1892) );
  XOR2_X1 U2172 ( .A(n2174), .B(n1892), .Z(mult_x_6_n1385) );
  AOI22_X1 U2173 ( .A1(mul_operand_b_q[27]), .A2(n2218), .B1(
        mul_operand_b_q[26]), .B2(n1020), .ZN(n1894) );
  AOI22_X1 U2174 ( .A1(mul_operand_b_q[25]), .A2(n2226), .B1(mult_x_6_n1077), 
        .B2(n2213), .ZN(n1893) );
  NAND2_X1 U2175 ( .A1(n1894), .A2(n1893), .ZN(n1895) );
  XOR2_X1 U2176 ( .A(n2174), .B(n1895), .Z(mult_x_6_n1386) );
  AOI22_X1 U2177 ( .A1(n2182), .A2(n2217), .B1(mul_operand_b_q[25]), .B2(n1020), .ZN(n1897) );
  AOI22_X1 U2178 ( .A1(n2183), .A2(n405), .B1(mult_x_6_n1078), .B2(n2213), 
        .ZN(n1896) );
  NAND2_X1 U2179 ( .A1(n1897), .A2(n1896), .ZN(n1898) );
  XOR2_X1 U2180 ( .A(n2174), .B(n1898), .Z(mult_x_6_n1387) );
  AOI22_X1 U2181 ( .A1(mul_operand_b_q[25]), .A2(n2218), .B1(
        mul_operand_b_q[24]), .B2(n2216), .ZN(n19001) );
  AOI22_X1 U2182 ( .A1(mul_operand_b_q[23]), .A2(n405), .B1(mult_x_6_n1079), 
        .B2(n2213), .ZN(n1899) );
  NAND2_X1 U2183 ( .A1(n19001), .A2(n1899), .ZN(n1901) );
  XOR2_X1 U2184 ( .A(n2174), .B(n1901), .Z(mult_x_6_n1388) );
  AOI22_X1 U2185 ( .A1(n2183), .A2(n2217), .B1(mul_operand_b_q[23]), .B2(n1020), .ZN(n1903) );
  AOI22_X1 U2186 ( .A1(mul_operand_b_q[22]), .A2(n2226), .B1(mult_x_6_n1080), 
        .B2(n2213), .ZN(n1902) );
  NAND2_X1 U2187 ( .A1(n1903), .A2(n1902), .ZN(n1904) );
  XOR2_X1 U2188 ( .A(n2174), .B(n1904), .Z(mult_x_6_n1389) );
  AOI22_X1 U2189 ( .A1(mul_operand_b_q[23]), .A2(n2218), .B1(
        mul_operand_b_q[22]), .B2(n1020), .ZN(n1906) );
  AOI22_X1 U2190 ( .A1(mul_operand_b_q[21]), .A2(n405), .B1(mult_x_6_n1081), 
        .B2(n2213), .ZN(n1905) );
  NAND2_X1 U2191 ( .A1(n1906), .A2(n1905), .ZN(n1907) );
  XOR2_X1 U2192 ( .A(n2174), .B(n1907), .Z(mult_x_6_n1390) );
  AOI22_X1 U2193 ( .A1(mul_operand_b_q[22]), .A2(n2217), .B1(
        mul_operand_b_q[21]), .B2(n1020), .ZN(n1909) );
  AOI22_X1 U2194 ( .A1(mul_operand_b_q[20]), .A2(n405), .B1(mult_x_6_n1082), 
        .B2(n2213), .ZN(n1908) );
  NAND2_X1 U2195 ( .A1(n1909), .A2(n1908), .ZN(n19101) );
  XOR2_X1 U2196 ( .A(n2174), .B(n19101), .Z(mult_x_6_n1391) );
  AOI22_X1 U2197 ( .A1(mul_operand_b_q[21]), .A2(n2218), .B1(
        mul_operand_b_q[20]), .B2(n1020), .ZN(n1912) );
  AOI22_X1 U2198 ( .A1(mul_operand_b_q[19]), .A2(n2226), .B1(mult_x_6_n1083), 
        .B2(n2213), .ZN(n1911) );
  NAND2_X1 U2199 ( .A1(n1912), .A2(n1911), .ZN(n1913) );
  XOR2_X1 U2200 ( .A(n2174), .B(n1913), .Z(mult_x_6_n1392) );
  AOI22_X1 U2201 ( .A1(mul_operand_b_q[20]), .A2(n2217), .B1(
        mul_operand_b_q[19]), .B2(n1020), .ZN(n1915) );
  AOI22_X1 U2202 ( .A1(mul_operand_b_q[18]), .A2(n405), .B1(mult_x_6_n1084), 
        .B2(n2213), .ZN(n1914) );
  NAND2_X1 U2203 ( .A1(n1915), .A2(n1914), .ZN(n1916) );
  XOR2_X1 U2204 ( .A(n2174), .B(n1916), .Z(mult_x_6_n1393) );
  AOI22_X1 U2205 ( .A1(mul_operand_b_q[19]), .A2(n2218), .B1(
        mul_operand_b_q[18]), .B2(n2216), .ZN(n1918) );
  AOI22_X1 U2206 ( .A1(mul_operand_b_q[17]), .A2(n405), .B1(mult_x_6_n1085), 
        .B2(n2213), .ZN(n1917) );
  NAND2_X1 U2207 ( .A1(n1918), .A2(n1917), .ZN(n1919) );
  XOR2_X1 U2208 ( .A(n2174), .B(n1919), .Z(mult_x_6_n1394) );
  AOI22_X1 U2209 ( .A1(mul_operand_b_q[17]), .A2(n1020), .B1(
        mul_operand_b_q[18]), .B2(n2217), .ZN(n1921) );
  AOI22_X1 U2210 ( .A1(n2185), .A2(n2226), .B1(mult_x_6_n1086), .B2(n2213), 
        .ZN(n19201) );
  NAND2_X1 U2211 ( .A1(n1921), .A2(n19201), .ZN(n1922) );
  XOR2_X1 U2212 ( .A(n2174), .B(n1922), .Z(mult_x_6_n1395) );
  AOI22_X1 U2213 ( .A1(mul_operand_b_q[17]), .A2(n2218), .B1(n2184), .B2(n1020), .ZN(n1924) );
  AOI22_X1 U2214 ( .A1(mul_operand_b_q[15]), .A2(n405), .B1(mult_x_6_n1087), 
        .B2(n2213), .ZN(n1923) );
  NAND2_X1 U2215 ( .A1(n1924), .A2(n1923), .ZN(n1925) );
  XOR2_X1 U2216 ( .A(n2174), .B(n1925), .Z(mult_x_6_n1396) );
  AOI22_X1 U2217 ( .A1(n2185), .A2(n2217), .B1(mul_operand_b_q[15]), .B2(n1020), .ZN(n1927) );
  AOI22_X1 U2218 ( .A1(mul_operand_b_q[14]), .A2(n405), .B1(mult_x_6_n1088), 
        .B2(n2213), .ZN(n1926) );
  NAND2_X1 U2219 ( .A1(n1927), .A2(n1926), .ZN(n1928) );
  XOR2_X1 U2220 ( .A(n2174), .B(n1928), .Z(mult_x_6_n1397) );
  AOI22_X1 U2221 ( .A1(mul_operand_b_q[15]), .A2(n2218), .B1(
        mul_operand_b_q[14]), .B2(n1020), .ZN(n19301) );
  AOI22_X1 U2222 ( .A1(mul_operand_b_q[13]), .A2(n2226), .B1(mult_x_6_n1089), 
        .B2(n2213), .ZN(n1929) );
  NAND2_X1 U2223 ( .A1(n19301), .A2(n1929), .ZN(n1931) );
  XOR2_X1 U2224 ( .A(n2174), .B(n1931), .Z(mult_x_6_n1398) );
  AOI22_X1 U2225 ( .A1(mul_operand_b_q[14]), .A2(n2218), .B1(
        mul_operand_b_q[13]), .B2(n1020), .ZN(n1933) );
  AOI22_X1 U2226 ( .A1(mul_operand_b_q[12]), .A2(n405), .B1(mult_x_6_n1090), 
        .B2(n2214), .ZN(n1932) );
  NAND2_X1 U2227 ( .A1(n1933), .A2(n1932), .ZN(n1934) );
  XOR2_X1 U2228 ( .A(n2174), .B(n1934), .Z(mult_x_6_n1399) );
  AOI22_X1 U2229 ( .A1(mul_operand_b_q[13]), .A2(n2217), .B1(
        mul_operand_b_q[12]), .B2(n1020), .ZN(n1936) );
  AOI22_X1 U2230 ( .A1(mul_operand_b_q[11]), .A2(n405), .B1(mult_x_6_n1091), 
        .B2(n2214), .ZN(n1935) );
  NAND2_X1 U2231 ( .A1(n1936), .A2(n1935), .ZN(n1937) );
  XOR2_X1 U2232 ( .A(n2174), .B(n1937), .Z(mult_x_6_n1400) );
  AOI22_X1 U2233 ( .A1(mul_operand_b_q[11]), .A2(n1020), .B1(
        mul_operand_b_q[12]), .B2(n2217), .ZN(n1939) );
  AOI22_X1 U2234 ( .A1(mul_operand_b_q[10]), .A2(n2226), .B1(mult_x_6_n1092), 
        .B2(n2214), .ZN(n1938) );
  NAND2_X1 U2235 ( .A1(n1939), .A2(n1938), .ZN(n19401) );
  XOR2_X1 U2236 ( .A(n2174), .B(n19401), .Z(mult_x_6_n1401) );
  AOI22_X1 U2237 ( .A1(mul_operand_b_q[11]), .A2(n2218), .B1(
        mul_operand_b_q[10]), .B2(n1020), .ZN(n1942) );
  AOI22_X1 U2238 ( .A1(n2187), .A2(n405), .B1(n2287), .B2(n2214), .ZN(n1941)
         );
  NAND2_X1 U2239 ( .A1(n1942), .A2(n1941), .ZN(n1943) );
  XOR2_X1 U2240 ( .A(n2174), .B(n1943), .Z(mult_x_6_n1402) );
  AOI22_X1 U2241 ( .A1(mul_operand_b_q[10]), .A2(n2217), .B1(n2186), .B2(n2216), .ZN(n1945) );
  AOI22_X1 U2242 ( .A1(mul_operand_b_q[8]), .A2(n405), .B1(mult_x_6_n1094), 
        .B2(n2213), .ZN(n1944) );
  NAND2_X1 U2243 ( .A1(n1945), .A2(n1944), .ZN(n1946) );
  XOR2_X1 U2244 ( .A(n2174), .B(n1946), .Z(mult_x_6_n1403) );
  AOI22_X1 U2245 ( .A1(n2187), .A2(n2218), .B1(mul_operand_b_q[8]), .B2(n1020), 
        .ZN(n1948) );
  AOI22_X1 U2246 ( .A1(mul_operand_b_q[7]), .A2(n2226), .B1(mult_x_6_n1095), 
        .B2(n2213), .ZN(n1947) );
  NAND2_X1 U2247 ( .A1(n1948), .A2(n1947), .ZN(n1949) );
  XOR2_X1 U2248 ( .A(n2174), .B(n1949), .Z(mult_x_6_n1404) );
  AOI22_X1 U2249 ( .A1(mul_operand_b_q[8]), .A2(n2217), .B1(mul_operand_b_q[7]), .B2(n1020), .ZN(n1951) );
  AOI22_X1 U2250 ( .A1(n2189), .A2(n405), .B1(mult_x_6_n1096), .B2(n2214), 
        .ZN(n19501) );
  NAND2_X1 U2251 ( .A1(n1951), .A2(n19501), .ZN(n1952) );
  XOR2_X1 U2252 ( .A(n2174), .B(n1952), .Z(mult_x_6_n1405) );
  AOI22_X1 U2253 ( .A1(mul_operand_b_q[7]), .A2(n2218), .B1(n2188), .B2(n1020), 
        .ZN(n1954) );
  AOI22_X1 U2254 ( .A1(n2190), .A2(n405), .B1(mult_x_6_n1097), .B2(n2214), 
        .ZN(n1953) );
  NAND2_X1 U2255 ( .A1(n1954), .A2(n1953), .ZN(n1955) );
  XOR2_X1 U2256 ( .A(n2174), .B(n1955), .Z(mult_x_6_n1406) );
  AOI22_X1 U2257 ( .A1(n2193), .A2(n2218), .B1(n1009), .B2(n1020), .ZN(n1957)
         );
  AOI22_X1 U2258 ( .A1(n2195), .A2(n2226), .B1(mult_x_6_n1101), .B2(n2214), 
        .ZN(n1956) );
  XOR2_X1 U2259 ( .A(mul_operand_a_q[5]), .B(mul_operand_a_q[4]), .Z(n1963) );
  XNOR2_X1 U2260 ( .A(mul_operand_a_q[4]), .B(mul_operand_a_q[3]), .ZN(n19601)
         );
  NAND2_X1 U2261 ( .A1(n1961), .A2(n2177), .ZN(n1962) );
  XOR2_X1 U2262 ( .A(n2175), .B(n1962), .Z(mult_x_6_n1414) );
  NOR2_X1 U2263 ( .A1(n2143), .A2(n1963), .ZN(n2048) );
  OR2_X1 U2264 ( .A1(n2223), .A2(n2221), .ZN(n1964) );
  AOI222_X1 U2265 ( .A1(n1964), .A2(mul_operand_b_q[32]), .B1(mult_x_6_n1071), 
        .B2(n2219), .C1(n2179), .C2(n624), .ZN(n1965) );
  XNOR2_X1 U2266 ( .A(n2175), .B(n1965), .ZN(mult_x_6_n1415) );
  AOI22_X1 U2267 ( .A1(n2180), .A2(n624), .B1(mult_x_6_n1072), .B2(n2219), 
        .ZN(n1967) );
  NAND2_X1 U2268 ( .A1(n2177), .A2(n2222), .ZN(n1966) );
  OAI211_X1 U2269 ( .C1(n2178), .C2(n2427), .A(n1967), .B(n1966), .ZN(n1968)
         );
  XOR2_X1 U2270 ( .A(n2175), .B(n1968), .Z(mult_x_6_n1416) );
  AOI22_X1 U2271 ( .A1(n2179), .A2(n2223), .B1(n2180), .B2(n2220), .ZN(n19701)
         );
  AOI22_X1 U2272 ( .A1(mul_operand_b_q[29]), .A2(n624), .B1(mult_x_6_n1073), 
        .B2(n2219), .ZN(n1969) );
  NAND2_X1 U2273 ( .A1(n19701), .A2(n1969), .ZN(n1971) );
  XOR2_X1 U2274 ( .A(n2175), .B(n1971), .Z(mult_x_6_n1417) );
  AOI22_X1 U2275 ( .A1(n2180), .A2(n2222), .B1(mul_operand_b_q[29]), .B2(n2221), .ZN(n1973) );
  AOI22_X1 U2276 ( .A1(n2181), .A2(n624), .B1(mult_x_6_n1074), .B2(n2219), 
        .ZN(n1972) );
  NAND2_X1 U2277 ( .A1(n1973), .A2(n1972), .ZN(n1974) );
  XOR2_X1 U2278 ( .A(n2175), .B(n1974), .Z(mult_x_6_n1418) );
  AOI22_X1 U2279 ( .A1(mul_operand_b_q[29]), .A2(n2223), .B1(
        mul_operand_b_q[28]), .B2(n2221), .ZN(n1976) );
  AOI22_X1 U2280 ( .A1(mul_operand_b_q[27]), .A2(n624), .B1(mult_x_6_n1075), 
        .B2(n2219), .ZN(n1975) );
  NAND2_X1 U2281 ( .A1(n1976), .A2(n1975), .ZN(n1977) );
  XOR2_X1 U2282 ( .A(n2175), .B(n1977), .Z(mult_x_6_n1419) );
  AOI22_X1 U2283 ( .A1(n2181), .A2(n2222), .B1(mul_operand_b_q[27]), .B2(n2221), .ZN(n1979) );
  AOI22_X1 U2284 ( .A1(n2182), .A2(n624), .B1(mult_x_6_n1076), .B2(n2219), 
        .ZN(n1978) );
  NAND2_X1 U2285 ( .A1(n1979), .A2(n1978), .ZN(n19801) );
  XOR2_X1 U2286 ( .A(n2175), .B(n19801), .Z(mult_x_6_n1420) );
  AOI22_X1 U2287 ( .A1(mul_operand_b_q[27]), .A2(n2223), .B1(
        mul_operand_b_q[26]), .B2(n2220), .ZN(n1982) );
  AOI22_X1 U2288 ( .A1(mul_operand_b_q[25]), .A2(n624), .B1(mult_x_6_n1077), 
        .B2(n2219), .ZN(n1981) );
  NAND2_X1 U2289 ( .A1(n1982), .A2(n1981), .ZN(n1983) );
  XOR2_X1 U2290 ( .A(n2175), .B(n1983), .Z(mult_x_6_n1421) );
  AOI22_X1 U2291 ( .A1(n2182), .A2(n2222), .B1(mul_operand_b_q[25]), .B2(n2221), .ZN(n1985) );
  AOI22_X1 U2292 ( .A1(n2183), .A2(n624), .B1(mult_x_6_n1078), .B2(n2219), 
        .ZN(n1984) );
  NAND2_X1 U2293 ( .A1(n1985), .A2(n1984), .ZN(n1986) );
  XOR2_X1 U2294 ( .A(n2175), .B(n1986), .Z(mult_x_6_n1422) );
  AOI22_X1 U2295 ( .A1(mul_operand_b_q[25]), .A2(n2223), .B1(
        mul_operand_b_q[24]), .B2(n2221), .ZN(n1988) );
  AOI22_X1 U2296 ( .A1(mul_operand_b_q[23]), .A2(n624), .B1(mult_x_6_n1079), 
        .B2(n2219), .ZN(n1987) );
  NAND2_X1 U2297 ( .A1(n1988), .A2(n1987), .ZN(n1989) );
  XOR2_X1 U2298 ( .A(n2175), .B(n1989), .Z(mult_x_6_n1423) );
  AOI22_X1 U2299 ( .A1(n2183), .A2(n2222), .B1(mul_operand_b_q[23]), .B2(n2221), .ZN(n1991) );
  AOI22_X1 U2300 ( .A1(mul_operand_b_q[22]), .A2(n624), .B1(mult_x_6_n1080), 
        .B2(n2219), .ZN(n19901) );
  NAND2_X1 U2301 ( .A1(n1991), .A2(n19901), .ZN(n1992) );
  XOR2_X1 U2302 ( .A(n2175), .B(n1992), .Z(mult_x_6_n1424) );
  AOI22_X1 U2303 ( .A1(mul_operand_b_q[23]), .A2(n2223), .B1(
        mul_operand_b_q[22]), .B2(n2220), .ZN(n1994) );
  AOI22_X1 U2304 ( .A1(mul_operand_b_q[21]), .A2(n624), .B1(mult_x_6_n1081), 
        .B2(n2219), .ZN(n1993) );
  NAND2_X1 U2305 ( .A1(n1994), .A2(n1993), .ZN(n1995) );
  XOR2_X1 U2306 ( .A(n2175), .B(n1995), .Z(mult_x_6_n1425) );
  AOI22_X1 U2307 ( .A1(mul_operand_b_q[22]), .A2(n2222), .B1(
        mul_operand_b_q[21]), .B2(n2221), .ZN(n1997) );
  AOI22_X1 U2308 ( .A1(mul_operand_b_q[20]), .A2(n624), .B1(mult_x_6_n1082), 
        .B2(n2219), .ZN(n1996) );
  NAND2_X1 U2309 ( .A1(n1997), .A2(n1996), .ZN(n1998) );
  XOR2_X1 U2310 ( .A(n2175), .B(n1998), .Z(mult_x_6_n1426) );
  AOI22_X1 U2311 ( .A1(mul_operand_b_q[21]), .A2(n2223), .B1(
        mul_operand_b_q[20]), .B2(n2221), .ZN(n20001) );
  AOI22_X1 U2312 ( .A1(mul_operand_b_q[19]), .A2(n624), .B1(mult_x_6_n1083), 
        .B2(n2219), .ZN(n1999) );
  NAND2_X1 U2313 ( .A1(n20001), .A2(n1999), .ZN(n2001) );
  XOR2_X1 U2314 ( .A(n2175), .B(n2001), .Z(mult_x_6_n1427) );
  AOI22_X1 U2315 ( .A1(mul_operand_b_q[20]), .A2(n2222), .B1(
        mul_operand_b_q[19]), .B2(n2221), .ZN(n2003) );
  AOI22_X1 U2316 ( .A1(mul_operand_b_q[18]), .A2(n624), .B1(mult_x_6_n1084), 
        .B2(n2219), .ZN(n2002) );
  NAND2_X1 U2317 ( .A1(n2003), .A2(n2002), .ZN(n2004) );
  XOR2_X1 U2318 ( .A(n2175), .B(n2004), .Z(mult_x_6_n1428) );
  AOI22_X1 U2319 ( .A1(mul_operand_b_q[19]), .A2(n2223), .B1(
        mul_operand_b_q[18]), .B2(n2220), .ZN(n2006) );
  AOI22_X1 U2320 ( .A1(mul_operand_b_q[17]), .A2(n624), .B1(mult_x_6_n1085), 
        .B2(n2219), .ZN(n2005) );
  NAND2_X1 U2321 ( .A1(n2006), .A2(n2005), .ZN(n2007) );
  XOR2_X1 U2322 ( .A(n2175), .B(n2007), .Z(mult_x_6_n1429) );
  AOI22_X1 U2323 ( .A1(mul_operand_b_q[17]), .A2(n2221), .B1(
        mul_operand_b_q[18]), .B2(n2222), .ZN(n2009) );
  AOI22_X1 U2324 ( .A1(n2185), .A2(n624), .B1(mult_x_6_n1086), .B2(n2219), 
        .ZN(n2008) );
  NAND2_X1 U2325 ( .A1(n2009), .A2(n2008), .ZN(n2010) );
  XOR2_X1 U2326 ( .A(n2175), .B(n2010), .Z(mult_x_6_n1430) );
  AOI22_X1 U2327 ( .A1(mul_operand_b_q[17]), .A2(n2223), .B1(n2184), .B2(n2221), .ZN(n2012) );
  AOI22_X1 U2328 ( .A1(mul_operand_b_q[15]), .A2(n624), .B1(mult_x_6_n1087), 
        .B2(n2219), .ZN(n2011) );
  NAND2_X1 U2329 ( .A1(n2012), .A2(n2011), .ZN(n2013) );
  XOR2_X1 U2330 ( .A(n2175), .B(n2013), .Z(mult_x_6_n1431) );
  AOI22_X1 U2331 ( .A1(n2185), .A2(n2223), .B1(mul_operand_b_q[15]), .B2(n2221), .ZN(n2015) );
  AOI22_X1 U2332 ( .A1(mul_operand_b_q[14]), .A2(n624), .B1(mult_x_6_n1088), 
        .B2(n2219), .ZN(n2014) );
  NAND2_X1 U2333 ( .A1(n2015), .A2(n2014), .ZN(n2016) );
  XOR2_X1 U2334 ( .A(n2176), .B(n2016), .Z(mult_x_6_n1432) );
  AOI22_X1 U2335 ( .A1(mul_operand_b_q[15]), .A2(n2222), .B1(
        mul_operand_b_q[14]), .B2(n2221), .ZN(n2018) );
  AOI22_X1 U2336 ( .A1(mul_operand_b_q[13]), .A2(n624), .B1(mult_x_6_n1089), 
        .B2(n2219), .ZN(n2017) );
  NAND2_X1 U2337 ( .A1(n2018), .A2(n2017), .ZN(n2019) );
  XOR2_X1 U2338 ( .A(n2176), .B(n2019), .Z(mult_x_6_n1433) );
  AOI22_X1 U2339 ( .A1(mul_operand_b_q[14]), .A2(n2223), .B1(
        mul_operand_b_q[13]), .B2(n2220), .ZN(n2021) );
  AOI22_X1 U2340 ( .A1(mul_operand_b_q[12]), .A2(n624), .B1(mult_x_6_n1090), 
        .B2(n2219), .ZN(n2020) );
  NAND2_X1 U2341 ( .A1(n2021), .A2(n2020), .ZN(n2022) );
  XOR2_X1 U2342 ( .A(n2176), .B(n2022), .Z(mult_x_6_n1434) );
  AOI22_X1 U2343 ( .A1(mul_operand_b_q[13]), .A2(n2222), .B1(
        mul_operand_b_q[12]), .B2(n2221), .ZN(n2024) );
  AOI22_X1 U2344 ( .A1(mul_operand_b_q[11]), .A2(n2144), .B1(mult_x_6_n1091), 
        .B2(n2219), .ZN(n2023) );
  NAND2_X1 U2345 ( .A1(n2024), .A2(n2023), .ZN(n2025) );
  XOR2_X1 U2346 ( .A(n2176), .B(n2025), .Z(mult_x_6_n1435) );
  AOI22_X1 U2347 ( .A1(mul_operand_b_q[11]), .A2(n2221), .B1(
        mul_operand_b_q[12]), .B2(n2222), .ZN(n2027) );
  AOI22_X1 U2348 ( .A1(mul_operand_b_q[10]), .A2(n2144), .B1(mult_x_6_n1092), 
        .B2(n2219), .ZN(n2026) );
  NAND2_X1 U2349 ( .A1(n2027), .A2(n2026), .ZN(n2028) );
  XOR2_X1 U2350 ( .A(n2176), .B(n2028), .Z(mult_x_6_n1436) );
  AOI22_X1 U2351 ( .A1(mul_operand_b_q[11]), .A2(n2222), .B1(
        mul_operand_b_q[10]), .B2(n2221), .ZN(n2030) );
  AOI22_X1 U2352 ( .A1(n2187), .A2(n2144), .B1(mult_x_6_n1093), .B2(n2219), 
        .ZN(n2029) );
  NAND2_X1 U2353 ( .A1(n2030), .A2(n2029), .ZN(n2031) );
  XOR2_X1 U2354 ( .A(n2176), .B(n2031), .Z(mult_x_6_n1437) );
  AOI22_X1 U2355 ( .A1(mul_operand_b_q[10]), .A2(n2223), .B1(n2186), .B2(n2221), .ZN(n2033) );
  AOI22_X1 U2356 ( .A1(mul_operand_b_q[8]), .A2(n2144), .B1(mult_x_6_n1094), 
        .B2(n2219), .ZN(n2032) );
  NAND2_X1 U2357 ( .A1(n2033), .A2(n2032), .ZN(n2034) );
  AOI22_X1 U2358 ( .A1(n2187), .A2(n2223), .B1(mul_operand_b_q[8]), .B2(n2221), 
        .ZN(n2036) );
  AOI22_X1 U2359 ( .A1(mul_operand_b_q[7]), .A2(n2144), .B1(mult_x_6_n1095), 
        .B2(n2219), .ZN(n2035) );
  NAND2_X1 U2360 ( .A1(n2036), .A2(n2035), .ZN(n2037) );
  XOR2_X1 U2361 ( .A(n2176), .B(n2037), .Z(mult_x_6_n1439) );
  AOI22_X1 U2362 ( .A1(mul_operand_b_q[8]), .A2(n2222), .B1(mul_operand_b_q[7]), .B2(n2221), .ZN(n2039) );
  AOI22_X1 U2363 ( .A1(n2189), .A2(n2144), .B1(mult_x_6_n1096), .B2(n2219), 
        .ZN(n2038) );
  NAND2_X1 U2364 ( .A1(n2039), .A2(n2038), .ZN(n2040) );
  XOR2_X1 U2365 ( .A(n2176), .B(n2040), .Z(mult_x_6_n1440) );
  AOI22_X1 U2366 ( .A1(mul_operand_b_q[7]), .A2(n2223), .B1(n2188), .B2(n2221), 
        .ZN(n2042) );
  AOI22_X1 U2367 ( .A1(n2190), .A2(n2144), .B1(mult_x_6_n1097), .B2(n2219), 
        .ZN(n2041) );
  NAND2_X1 U2368 ( .A1(n2042), .A2(n2041), .ZN(n2043) );
  XOR2_X1 U2369 ( .A(n2175), .B(n2043), .Z(mult_x_6_n1441) );
  AOI22_X1 U2370 ( .A1(n2193), .A2(n2223), .B1(n1009), .B2(n2220), .ZN(n2044)
         );
  XOR2_X1 U2371 ( .A(n2176), .B(n2045), .Z(mult_x_6_n1445) );
  AOI22_X1 U2372 ( .A1(n1009), .A2(n2048), .B1(n2286), .B2(n2220), .ZN(n2046)
         );
  NOR3_X1 U2373 ( .A1(mul_operand_a_q[1]), .A2(mul_operand_a_q[0]), .A3(n1025), 
        .ZN(n2119) );
  AOI22_X1 U2374 ( .A1(n2179), .A2(n385), .B1(n2180), .B2(n608), .ZN(n2051) );
  AOI22_X1 U2375 ( .A1(n2225), .A2(mult_x_6_n1073), .B1(n2224), .B2(
        mul_operand_b_q[29]), .ZN(n2050) );
  NAND2_X1 U2376 ( .A1(n2051), .A2(n2050), .ZN(n2052) );
  XNOR2_X1 U2377 ( .A(n2052), .B(n1013), .ZN(mult_x_6_n1452) );
  AOI22_X1 U2378 ( .A1(n2180), .A2(n385), .B1(n608), .B2(mul_operand_b_q[29]), 
        .ZN(n2054) );
  AOI22_X1 U2379 ( .A1(n2225), .A2(mult_x_6_n1074), .B1(n2224), .B2(
        mul_operand_b_q[28]), .ZN(n2053) );
  NAND2_X1 U2380 ( .A1(n2054), .A2(n2053), .ZN(n2055) );
  AOI22_X1 U2381 ( .A1(n385), .A2(mul_operand_b_q[29]), .B1(n608), .B2(
        mul_operand_b_q[28]), .ZN(n2057) );
  AOI22_X1 U2382 ( .A1(n2225), .A2(mult_x_6_n1075), .B1(n2224), .B2(
        mul_operand_b_q[27]), .ZN(n2056) );
  NAND2_X1 U2383 ( .A1(n2057), .A2(n2056), .ZN(n2058) );
  XNOR2_X1 U2384 ( .A(n2058), .B(n1013), .ZN(mult_x_6_n1454) );
  AOI22_X1 U2385 ( .A1(n385), .A2(mul_operand_b_q[28]), .B1(n608), .B2(
        mul_operand_b_q[27]), .ZN(n2060) );
  AOI22_X1 U2386 ( .A1(n2225), .A2(mult_x_6_n1076), .B1(n2224), .B2(
        mul_operand_b_q[26]), .ZN(n2059) );
  NAND2_X1 U2387 ( .A1(n2060), .A2(n2059), .ZN(n2061) );
  XNOR2_X1 U2388 ( .A(n2061), .B(n1013), .ZN(mult_x_6_n1455) );
  AOI22_X1 U2389 ( .A1(n385), .A2(mul_operand_b_q[27]), .B1(n608), .B2(
        mul_operand_b_q[26]), .ZN(n2063) );
  AOI22_X1 U2390 ( .A1(n2225), .A2(mult_x_6_n1077), .B1(n2224), .B2(
        mul_operand_b_q[25]), .ZN(n2062) );
  NAND2_X1 U2391 ( .A1(n2063), .A2(n2062), .ZN(n2064) );
  AOI22_X1 U2392 ( .A1(n385), .A2(mul_operand_b_q[25]), .B1(n608), .B2(n2183), 
        .ZN(n2066) );
  AOI22_X1 U2393 ( .A1(n2225), .A2(mult_x_6_n1079), .B1(n2224), .B2(
        mul_operand_b_q[23]), .ZN(n2065) );
  NAND2_X1 U2394 ( .A1(n2066), .A2(n2065), .ZN(n2067) );
  XNOR2_X1 U2395 ( .A(n2067), .B(n1013), .ZN(mult_x_6_n1458) );
  AOI22_X1 U2396 ( .A1(n385), .A2(n2183), .B1(n608), .B2(mul_operand_b_q[23]), 
        .ZN(n2069) );
  AOI22_X1 U2397 ( .A1(n2225), .A2(mult_x_6_n1080), .B1(n2224), .B2(
        mul_operand_b_q[22]), .ZN(n2068) );
  NAND2_X1 U2398 ( .A1(n2069), .A2(n2068), .ZN(n2070) );
  XNOR2_X1 U2399 ( .A(n2070), .B(n1013), .ZN(mult_x_6_n1459) );
  AOI22_X1 U2400 ( .A1(n385), .A2(mul_operand_b_q[23]), .B1(n608), .B2(
        mul_operand_b_q[22]), .ZN(n2072) );
  AOI22_X1 U2401 ( .A1(n2225), .A2(mult_x_6_n1081), .B1(n2224), .B2(
        mul_operand_b_q[21]), .ZN(n2071) );
  NAND2_X1 U2402 ( .A1(n2072), .A2(n2071), .ZN(n2073) );
  XNOR2_X1 U2403 ( .A(n2073), .B(n1013), .ZN(mult_x_6_n1460) );
  AOI22_X1 U2404 ( .A1(n385), .A2(mul_operand_b_q[22]), .B1(n608), .B2(
        mul_operand_b_q[21]), .ZN(n2075) );
  AOI22_X1 U2405 ( .A1(n2225), .A2(mult_x_6_n1082), .B1(n2224), .B2(
        mul_operand_b_q[20]), .ZN(n2074) );
  NAND2_X1 U2406 ( .A1(n2075), .A2(n2074), .ZN(n2076) );
  XNOR2_X1 U2407 ( .A(n2076), .B(n1013), .ZN(mult_x_6_n1461) );
  AOI22_X1 U2408 ( .A1(n385), .A2(mul_operand_b_q[21]), .B1(n608), .B2(
        mul_operand_b_q[20]), .ZN(n2078) );
  AOI22_X1 U2409 ( .A1(n2225), .A2(mult_x_6_n1083), .B1(n2224), .B2(
        mul_operand_b_q[19]), .ZN(n2077) );
  NAND2_X1 U2410 ( .A1(n2078), .A2(n2077), .ZN(n2079) );
  XNOR2_X1 U2411 ( .A(n2079), .B(n1013), .ZN(mult_x_6_n1462) );
  AOI22_X1 U2412 ( .A1(n385), .A2(mul_operand_b_q[20]), .B1(n608), .B2(
        mul_operand_b_q[19]), .ZN(n2081) );
  AOI22_X1 U2413 ( .A1(n2225), .A2(mult_x_6_n1084), .B1(n2224), .B2(
        mul_operand_b_q[18]), .ZN(n2080) );
  NAND2_X1 U2414 ( .A1(n2081), .A2(n2080), .ZN(n2082) );
  XNOR2_X1 U2415 ( .A(n2082), .B(n1013), .ZN(mult_x_6_n1463) );
  AOI22_X1 U2416 ( .A1(n385), .A2(mul_operand_b_q[19]), .B1(n608), .B2(
        mul_operand_b_q[18]), .ZN(n2084) );
  AOI22_X1 U2417 ( .A1(n2225), .A2(mult_x_6_n1085), .B1(n2224), .B2(
        mul_operand_b_q[17]), .ZN(n2083) );
  NAND2_X1 U2418 ( .A1(n2084), .A2(n2083), .ZN(n2085) );
  XNOR2_X1 U2419 ( .A(n2085), .B(n1013), .ZN(mult_x_6_n1464) );
  AOI22_X1 U2420 ( .A1(n385), .A2(mul_operand_b_q[18]), .B1(n608), .B2(
        mul_operand_b_q[17]), .ZN(n2087) );
  AOI22_X1 U2421 ( .A1(n2225), .A2(mult_x_6_n1086), .B1(n2224), .B2(n2184), 
        .ZN(n2086) );
  NAND2_X1 U2422 ( .A1(n2087), .A2(n2086), .ZN(n2088) );
  XNOR2_X1 U2423 ( .A(n2088), .B(n1013), .ZN(mult_x_6_n1465) );
  AOI22_X1 U2424 ( .A1(n385), .A2(mul_operand_b_q[17]), .B1(n608), .B2(n2184), 
        .ZN(n2090) );
  AOI22_X1 U2425 ( .A1(n2225), .A2(mult_x_6_n1087), .B1(n2224), .B2(
        mul_operand_b_q[15]), .ZN(n2089) );
  NAND2_X1 U2426 ( .A1(n2090), .A2(n2089), .ZN(n2091) );
  XNOR2_X1 U2427 ( .A(n2091), .B(n1013), .ZN(mult_x_6_n1466) );
  AOI22_X1 U2428 ( .A1(n385), .A2(n2184), .B1(n608), .B2(mul_operand_b_q[15]), 
        .ZN(n2093) );
  AOI22_X1 U2429 ( .A1(n2225), .A2(mult_x_6_n1088), .B1(n2224), .B2(
        mul_operand_b_q[14]), .ZN(n2092) );
  NAND2_X1 U2430 ( .A1(n2092), .A2(n2093), .ZN(n2094) );
  XNOR2_X1 U2431 ( .A(n2094), .B(n1013), .ZN(mult_x_6_n1467) );
  AOI22_X1 U2432 ( .A1(n385), .A2(mul_operand_b_q[15]), .B1(n608), .B2(
        mul_operand_b_q[14]), .ZN(n2096) );
  AOI22_X1 U2433 ( .A1(n2225), .A2(mult_x_6_n1089), .B1(n2224), .B2(
        mul_operand_b_q[13]), .ZN(n2095) );
  NAND2_X1 U2434 ( .A1(n2096), .A2(n2095), .ZN(n2097) );
  XNOR2_X1 U2435 ( .A(n2097), .B(n1013), .ZN(mult_x_6_n1468) );
  AOI22_X1 U2436 ( .A1(n385), .A2(mul_operand_b_q[14]), .B1(n608), .B2(
        mul_operand_b_q[13]), .ZN(n2099) );
  AOI22_X1 U2437 ( .A1(n2225), .A2(mult_x_6_n1090), .B1(n2224), .B2(
        mul_operand_b_q[12]), .ZN(n2098) );
  NAND2_X1 U2438 ( .A1(n2099), .A2(n2098), .ZN(n2100) );
  XNOR2_X1 U2439 ( .A(n2100), .B(n1013), .ZN(mult_x_6_n1469) );
  AOI22_X1 U2440 ( .A1(n385), .A2(mul_operand_b_q[13]), .B1(n608), .B2(
        mul_operand_b_q[12]), .ZN(n2102) );
  AOI22_X1 U2441 ( .A1(n2225), .A2(mult_x_6_n1091), .B1(n2224), .B2(
        mul_operand_b_q[11]), .ZN(n2101) );
  NAND2_X1 U2442 ( .A1(n2102), .A2(n2101), .ZN(n2103) );
  XNOR2_X1 U2443 ( .A(n2103), .B(n1013), .ZN(mult_x_6_n1470) );
  AOI22_X1 U2444 ( .A1(n385), .A2(mul_operand_b_q[12]), .B1(n608), .B2(
        mul_operand_b_q[11]), .ZN(n2105) );
  AOI22_X1 U2445 ( .A1(n2225), .A2(mult_x_6_n1092), .B1(n2224), .B2(
        mul_operand_b_q[10]), .ZN(n2104) );
  NAND2_X1 U2446 ( .A1(n2105), .A2(n2104), .ZN(n2106) );
  XNOR2_X1 U2447 ( .A(n2106), .B(n1013), .ZN(mult_x_6_n1471) );
  AOI22_X1 U2448 ( .A1(n385), .A2(mul_operand_b_q[11]), .B1(n608), .B2(
        mul_operand_b_q[10]), .ZN(n2108) );
  AOI22_X1 U2449 ( .A1(n2225), .A2(mult_x_6_n1093), .B1(n2224), .B2(n2186), 
        .ZN(n2107) );
  NAND2_X1 U2450 ( .A1(n2108), .A2(n2107), .ZN(n2109) );
  XNOR2_X1 U2451 ( .A(n2109), .B(n1013), .ZN(mult_x_6_n1472) );
  AOI22_X1 U2452 ( .A1(n385), .A2(mul_operand_b_q[10]), .B1(n608), .B2(n2186), 
        .ZN(n2111) );
  AOI22_X1 U2453 ( .A1(n2225), .A2(mult_x_6_n1094), .B1(n2224), .B2(
        mul_operand_b_q[8]), .ZN(n2110) );
  NAND2_X1 U2454 ( .A1(n2111), .A2(n2110), .ZN(n2112) );
  XNOR2_X1 U2455 ( .A(n2112), .B(n1013), .ZN(mult_x_6_n1473) );
  AOI22_X1 U2456 ( .A1(n385), .A2(mul_operand_b_q[7]), .B1(n608), .B2(n2189), 
        .ZN(n2114) );
  AOI22_X1 U2457 ( .A1(mult_x_6_n1097), .A2(n2225), .B1(n2224), .B2(n2190), 
        .ZN(n2113) );
  NAND2_X1 U2458 ( .A1(n2114), .A2(n2113), .ZN(n2115) );
  XNOR2_X1 U2459 ( .A(n2115), .B(n1013), .ZN(mult_x_6_n1476) );
  AOI22_X1 U2460 ( .A1(n385), .A2(n2190), .B1(n608), .B2(n2192), .ZN(n2116) );
  AOI22_X1 U2461 ( .A1(n385), .A2(n2192), .B1(n608), .B2(n2193), .ZN(n2117) );
  XNOR2_X1 U2462 ( .A(n2118), .B(n1013), .ZN(mult_x_6_n1479) );
  AOI222_X1 U2463 ( .A1(n2120), .A2(mult_x_6_n1103), .B1(n2142), .B2(n2286), 
        .C1(n2141), .C2(n2196), .ZN(n2121) );
  XNOR2_X1 U2464 ( .A(n2122), .B(mul_operand_a_q[32]), .ZN(mult_x_6_n333) );
  AOI22_X1 U2465 ( .A1(n604), .A2(mul_operand_b_q[26]), .B1(n632), .B2(
        mul_operand_b_q[25]), .ZN(n2124) );
  AOI22_X1 U2466 ( .A1(n2132), .A2(mul_operand_b_q[24]), .B1(n2134), .B2(
        mult_x_6_n1078), .ZN(n2123) );
  NAND2_X1 U2467 ( .A1(n2124), .A2(n2123), .ZN(n2125) );
  XOR2_X1 U2468 ( .A(mul_operand_a_q[32]), .B(n2125), .Z(mult_x_6_n350) );
  AOI22_X1 U2469 ( .A1(n604), .A2(mul_operand_b_q[20]), .B1(n2132), .B2(
        mul_operand_b_q[18]), .ZN(n2127) );
  AOI22_X1 U2470 ( .A1(n632), .A2(mul_operand_b_q[19]), .B1(n2134), .B2(
        mult_x_6_n1084), .ZN(n2126) );
  NAND2_X1 U2471 ( .A1(n2127), .A2(n2126), .ZN(n2128) );
  XOR2_X1 U2472 ( .A(mul_operand_a_q[32]), .B(n2128), .Z(mult_x_6_n393) );
  AOI22_X1 U2473 ( .A1(n604), .A2(mul_operand_b_q[14]), .B1(n2132), .B2(
        mul_operand_b_q[12]), .ZN(n2130) );
  AOI22_X1 U2474 ( .A1(n632), .A2(mul_operand_b_q[13]), .B1(n2134), .B2(
        mult_x_6_n1090), .ZN(n2129) );
  NAND2_X1 U2475 ( .A1(n2130), .A2(n2129), .ZN(n2131) );
  XOR2_X1 U2476 ( .A(mul_operand_a_q[32]), .B(n2131), .Z(mult_x_6_n460) );
  AOI22_X1 U2477 ( .A1(n604), .A2(mul_operand_b_q[8]), .B1(n2132), .B2(n2189), 
        .ZN(n2137) );
  AOI22_X1 U2478 ( .A1(n632), .A2(mul_operand_b_q[7]), .B1(n2134), .B2(
        mult_x_6_n1096), .ZN(n2136) );
  NAND2_X1 U2479 ( .A1(n2137), .A2(n2136), .ZN(n2138) );
  XOR2_X1 U2480 ( .A(mul_operand_a_q[32]), .B(n2138), .Z(mult_x_6_n551) );
  OAI211_X1 U2481 ( .C1(mul_operand_a_q[1]), .C2(mul_operand_a_q[0]), .A(n2177), .B(n1013), .ZN(n2139) );
  OAI21_X1 U2482 ( .B1(n2177), .B2(n1013), .A(n2139), .ZN(n2140) );
  NAND2_X1 U2483 ( .A1(n2164), .A2(n2140), .ZN(mult_x_6_n606) );
  XOR2_X1 U2484 ( .A(mult_x_6_n664), .B(n2140), .Z(mult_x_6_n645) );
  INV_X1 U2485 ( .A(n2417), .ZN(n2198) );
  INV_X1 U2486 ( .A(n2426), .ZN(n2205) );
  INV_X1 U2487 ( .A(n2215), .ZN(n2216) );
  INV_X1 U2488 ( .A(n2427), .ZN(n2220) );
  NAND2_X1 U2489 ( .A1(mult_x_6_n1473), .A2(mult_x_6_n967), .ZN(n2227) );
  XOR2_X1 U2490 ( .A(mult_x_6_n321), .B(n2228), .Z(mult_result_w[10]) );
  XOR2_X1 U2491 ( .A(mult_x_6_n1473), .B(mult_x_6_n967), .Z(n2228) );
  NAND2_X1 U2492 ( .A1(mult_x_6_n1459), .A2(mult_x_6_n813), .ZN(n2229) );
  XOR2_X1 U2493 ( .A(mult_x_6_n307), .B(n2230), .Z(mult_result_w[24]) );
  XOR2_X1 U2494 ( .A(mult_x_6_n1459), .B(mult_x_6_n813), .Z(n2230) );
  XOR2_X1 U2495 ( .A(n1016), .B(n2231), .Z(mult_result_w[38]) );
  XOR2_X1 U2496 ( .A(mult_x_6_n554), .B(mult_x_6_n570), .Z(n2231) );
  XOR2_X1 U2497 ( .A(mult_x_6_n280), .B(n2232), .Z(mult_result_w[51]) );
  XOR2_X1 U2498 ( .A(mult_x_6_n386), .B(mult_x_6_n395), .Z(n2232) );
  NAND2_X1 U2499 ( .A1(n2187), .A2(mul_operand_b_q[10]), .ZN(n2233) );
  NAND3_X1 U2500 ( .A1(n2236), .A2(n2235), .A3(n2234), .ZN(mult_x_6_n1047) );
  NAND2_X1 U2501 ( .A1(mul_operand_b_q[23]), .A2(n2183), .ZN(n2234) );
  NAND2_X1 U2502 ( .A1(n2250), .A2(n2183), .ZN(n2235) );
  XOR2_X1 U2503 ( .A(n2250), .B(n2237), .Z(mult_x_6_n1080) );
  XOR2_X1 U2504 ( .A(mul_operand_b_q[23]), .B(n2183), .Z(n2237) );
  NAND2_X1 U2505 ( .A1(mult_x_6_n1451), .A2(mult_x_6_n667), .ZN(n2238) );
  XOR2_X1 U2506 ( .A(mult_x_6_n285), .B(n2239), .Z(mult_result_w[46]) );
  XOR2_X1 U2507 ( .A(mult_x_6_n448), .B(mult_x_6_n438), .Z(n2239) );
  NAND2_X1 U2508 ( .A1(mult_x_6_n336), .A2(mult_x_6_n335), .ZN(n2240) );
  XOR2_X1 U2509 ( .A(mult_x_6_n336), .B(mult_x_6_n335), .Z(n2241) );
  XOR2_X1 U2510 ( .A(mult_x_6_n333), .B(mult_x_6_n334), .Z(n2242) );
  XOR2_X1 U2511 ( .A(mult_x_6_n286), .B(n2243), .Z(mult_result_w[45]) );
  XOR2_X1 U2512 ( .A(mult_x_6_n449), .B(mult_x_6_n462), .Z(n2243) );
  NAND2_X1 U2513 ( .A1(n2187), .A2(mul_operand_b_q[8]), .ZN(n2244) );
  XOR2_X1 U2514 ( .A(n2187), .B(mul_operand_b_q[8]), .Z(n2247) );
  XOR2_X1 U2515 ( .A(mult_x_6_n1049), .B(n2248), .Z(mult_x_6_n1081) );
  XOR2_X1 U2516 ( .A(mul_operand_b_q[23]), .B(mul_operand_b_q[22]), .Z(n2248)
         );
  XOR2_X1 U2517 ( .A(n641), .B(n2249), .Z(mult_result_w[42]) );
  XOR2_X1 U2518 ( .A(mult_x_6_n490), .B(mult_x_6_n505), .Z(n2249) );
  NAND2_X1 U2519 ( .A1(mul_operand_b_q[8]), .A2(mul_operand_b_q[7]), .ZN(n2251) );
  XOR2_X1 U2520 ( .A(mult_x_6_n1053), .B(n2255), .Z(mult_x_6_n1085) );
  XOR2_X1 U2521 ( .A(mul_operand_b_q[19]), .B(mul_operand_b_q[18]), .Z(n2255)
         );
  XOR2_X1 U2522 ( .A(mult_x_6_n1042), .B(n2256), .Z(mult_x_6_n1074) );
  XOR2_X1 U2523 ( .A(mul_operand_b_q[29]), .B(mul_operand_b_q[30]), .Z(n2256)
         );
  NAND2_X1 U2524 ( .A1(n1009), .A2(n2194), .ZN(n2257) );
  NAND2_X1 U2525 ( .A1(mult_x_6_n1069), .A2(n2194), .ZN(n2258) );
  NAND2_X1 U2526 ( .A1(mult_x_6_n1069), .A2(n1009), .ZN(n2259) );
  NAND2_X1 U2527 ( .A1(mult_x_6_n1458), .A2(mult_x_6_n797), .ZN(n2260) );
  XOR2_X1 U2528 ( .A(mult_x_6_n306), .B(n2261), .Z(mult_result_w[25]) );
  XOR2_X1 U2529 ( .A(mult_x_6_n1458), .B(mult_x_6_n797), .Z(n2261) );
  NAND2_X1 U2530 ( .A1(mult_x_6_n1453), .A2(mult_x_6_n707), .ZN(n2262) );
  XOR2_X1 U2531 ( .A(mult_x_6_n275), .B(n2263), .Z(mult_result_w[56]) );
  XOR2_X1 U2532 ( .A(mult_x_6_n353), .B(mult_x_6_n357), .Z(n2263) );
  XOR2_X1 U2533 ( .A(mult_x_6_n1055), .B(n2264), .Z(mult_x_6_n1087) );
  XOR2_X1 U2534 ( .A(n2185), .B(mul_operand_b_q[17]), .Z(n2264) );
  NAND3_X1 U2535 ( .A1(n2267), .A2(n2266), .A3(n2265), .ZN(mult_x_6_n1040) );
  NAND2_X1 U2536 ( .A1(n2179), .A2(n2180), .ZN(n2265) );
  NAND2_X1 U2537 ( .A1(mult_x_6_n1041), .A2(n2180), .ZN(n2266) );
  NAND2_X1 U2538 ( .A1(mult_x_6_n1041), .A2(n2179), .ZN(n2267) );
  XOR2_X1 U2539 ( .A(n2179), .B(mul_operand_b_q[30]), .Z(n2268) );
  XOR2_X1 U2540 ( .A(mult_x_6_n277), .B(n2269), .Z(mult_result_w[54]) );
  XOR2_X1 U2541 ( .A(mult_x_6_n364), .B(mult_x_6_n371), .Z(n2269) );
  NAND2_X1 U2542 ( .A1(mult_x_6_n1471), .A2(mult_x_6_n953), .ZN(n2270) );
  XOR2_X1 U2543 ( .A(n1012), .B(n2271), .Z(mult_result_w[35]) );
  XOR2_X1 U2544 ( .A(mult_x_6_n609), .B(mult_x_6_n627), .Z(n2271) );
  NAND2_X1 U2545 ( .A1(mult_x_6_n1468), .A2(mult_x_6_n927), .ZN(n2272) );
  NAND2_X1 U2546 ( .A1(mult_x_6_n1463), .A2(mult_x_6_n871), .ZN(n2273) );
  XOR2_X1 U2547 ( .A(n1011), .B(n2274), .Z(mult_result_w[20]) );
  XOR2_X1 U2548 ( .A(mult_x_6_n1463), .B(mult_x_6_n871), .Z(n2274) );
  XOR2_X1 U2549 ( .A(mult_x_6_n1044), .B(n2276), .Z(mult_x_6_n1076) );
  XOR2_X1 U2550 ( .A(mul_operand_b_q[27]), .B(n2181), .Z(n2276) );
  NAND2_X1 U2551 ( .A1(mul_operand_b_q[25]), .A2(n2182), .ZN(n2277) );
  NAND2_X1 U2552 ( .A1(mult_x_6_n1046), .A2(n2182), .ZN(n2278) );
  NAND2_X1 U2553 ( .A1(mult_x_6_n1046), .A2(mul_operand_b_q[25]), .ZN(n2279)
         );
  XOR2_X1 U2554 ( .A(mult_x_6_n1046), .B(n2280), .Z(mult_x_6_n1078) );
  XOR2_X1 U2555 ( .A(mul_operand_b_q[25]), .B(n2182), .Z(n2280) );
  NAND2_X1 U2556 ( .A1(n2191), .A2(n2189), .ZN(n2281) );
  NAND2_X1 U2557 ( .A1(n2192), .A2(n2191), .ZN(n2282) );
  XOR2_X1 U2558 ( .A(mul_operand_b_q[4]), .B(n2191), .Z(n2285) );
  INV_X1 U2559 ( .A(n2242), .ZN(n2309) );
  INV_X1 U2560 ( .A(mult_x_6_n321), .ZN(n2314) );
  NOR2_X1 U2561 ( .A1(mult_x_6_n1473), .A2(mult_x_6_n967), .ZN(n2315) );
  NAND4_X1 U2562 ( .A1(n2246), .A2(n2245), .A3(n2319), .A4(n2322), .ZN(n2325)
         );
  XNOR2_X1 U2563 ( .A(mult_x_6_n856), .B(n2326), .ZN(mult_x_6_n843) );
  OR2_X1 U2564 ( .A1(mult_x_6_n813), .A2(mult_x_6_n1459), .ZN(n2328) );
  XNOR2_X1 U2565 ( .A(mult_x_6_n870), .B(n2330), .ZN(mult_x_6_n857) );
  OAI21_X1 U2566 ( .B1(n2341), .B2(n2340), .A(n2270), .ZN(mult_x_6_n318) );
  XNOR2_X1 U2567 ( .A(mult_x_6_n686), .B(n2344), .ZN(mult_x_6_n667) );
  NAND2_X1 U2568 ( .A1(mult_x_6_n669), .A2(mult_x_6_n1419), .ZN(n2346) );
  NAND2_X1 U2569 ( .A1(n2345), .A2(n2346), .ZN(mult_x_6_n666) );
  NAND2_X1 U2570 ( .A1(mult_x_6_n307), .A2(n2328), .ZN(n2347) );
  NAND2_X1 U2571 ( .A1(n2347), .A2(n2229), .ZN(mult_x_6_n306) );
  OAI21_X1 U2572 ( .B1(mult_x_6_n797), .B2(mult_x_6_n1458), .A(mult_x_6_n306), 
        .ZN(n2348) );
  XNOR2_X1 U2573 ( .A(mult_x_6_n812), .B(n2349), .ZN(mult_x_6_n797) );
  OR2_X1 U2574 ( .A1(mult_x_6_n799), .A2(mult_x_6_n1426), .ZN(n2350) );
  NAND2_X1 U2575 ( .A1(mult_x_6_n812), .A2(n2350), .ZN(n2351) );
  NAND2_X1 U2576 ( .A1(mult_x_6_n1475), .A2(mult_x_6_n979), .ZN(n2353) );
  XNOR2_X1 U2577 ( .A(n2359), .B(mult_x_6_n947), .ZN(n2354) );
  XNOR2_X1 U2578 ( .A(n2357), .B(n2358), .ZN(mult_x_6_n937) );
  INV_X1 U2579 ( .A(mult_x_6_n316), .ZN(n2361) );
  NOR2_X1 U2580 ( .A1(mult_x_6_n1468), .A2(mult_x_6_n927), .ZN(n2362) );
  XNOR2_X1 U2581 ( .A(mult_x_6_n688), .B(n2363), .ZN(mult_x_6_n669) );
  INV_X1 U2582 ( .A(mult_x_6_n299), .ZN(n2373) );
  NOR2_X1 U2583 ( .A1(mult_x_6_n667), .A2(mult_x_6_n1451), .ZN(n2374) );
  NOR2_X1 U2584 ( .A1(mult_x_6_n871), .A2(mult_x_6_n1463), .ZN(n2376) );
  NOR2_X1 U2585 ( .A1(mult_x_6_n651), .A2(mult_x_6_n1386), .ZN(n2380) );
  NAND2_X1 U2586 ( .A1(mult_x_6_n651), .A2(mult_x_6_n1386), .ZN(n2381) );
  OAI21_X1 U2587 ( .B1(n2380), .B2(n2379), .A(n2381), .ZN(mult_x_6_n648) );
  OR2_X1 U2588 ( .A1(mult_x_6_n845), .A2(mult_x_6_n1429), .ZN(n2382) );
  XNOR2_X1 U2589 ( .A(n2383), .B(mult_x_6_n746), .ZN(mult_x_6_n729) );
  INV_X1 U2590 ( .A(mult_x_6_n746), .ZN(n2385) );
  OAI21_X1 U2591 ( .B1(n2385), .B2(n2421), .A(n2384), .ZN(mult_x_6_n728) );
  NAND4_X1 U2592 ( .A1(n2283), .A2(n2284), .A3(n2389), .A4(n2392), .ZN(n2393)
         );
  NAND2_X1 U2593 ( .A1(n2391), .A2(n2388), .ZN(n2394) );
  NAND2_X1 U2594 ( .A1(n2394), .A2(n2389), .ZN(n2395) );
  NAND2_X1 U2595 ( .A1(mult_x_6_n323), .A2(n2398), .ZN(n2352) );
  XNOR2_X1 U2596 ( .A(mult_x_6_n946), .B(n2400), .ZN(mult_x_6_n939) );
  XNOR2_X1 U2597 ( .A(mult_x_6_n982), .B(n2402), .ZN(mult_x_6_n979) );
  NAND2_X1 U2598 ( .A1(mult_x_6_n982), .A2(n2424), .ZN(n2404) );
  NAND2_X1 U2599 ( .A1(n2404), .A2(n2403), .ZN(mult_x_6_n978) );
  NAND2_X1 U2600 ( .A1(n2407), .A2(n2262), .ZN(mult_x_6_n300) );
  OAI21_X1 U2601 ( .B1(mult_x_6_n707), .B2(mult_x_6_n1453), .A(mult_x_6_n301), 
        .ZN(n2407) );
  NAND2_X1 U2602 ( .A1(mult_x_6_n535), .A2(mult_x_6_n521), .ZN(n2408) );
  NAND2_X1 U2603 ( .A1(mult_x_6_n364), .A2(mult_x_6_n371), .ZN(n2409) );
  NAND2_X1 U2604 ( .A1(mult_x_6_n554), .A2(mult_x_6_n570), .ZN(n2410) );
  NAND2_X1 U2605 ( .A1(mult_x_6_n386), .A2(mult_x_6_n395), .ZN(n2411) );
  NAND2_X1 U2606 ( .A1(mult_x_6_n353), .A2(mult_x_6_n357), .ZN(n2412) );
  NAND2_X1 U2607 ( .A1(mult_x_6_n490), .A2(mult_x_6_n505), .ZN(n2413) );
  INV_X1 U2608 ( .A(n2288), .ZN(n2289) );
  INV_X1 U2609 ( .A(n2429), .ZN(n2365) );
  NAND2_X1 U2610 ( .A1(mult_x_6_n609), .A2(mult_x_6_n627), .ZN(n2420) );
  NOR2_X1 U2611 ( .A1(mult_x_6_n731), .A2(mult_x_6_n1390), .ZN(n2421) );
  NOR2_X1 U2612 ( .A1(mult_x_6_n817), .A2(mult_x_6_n1395), .ZN(n2422) );
  NAND2_X1 U2613 ( .A1(mult_x_6_n799), .A2(mult_x_6_n1426), .ZN(n2423) );
  OR2_X1 U2614 ( .A1(mult_x_6_n1443), .A2(mult_x_6_n981), .ZN(n2424) );
  INV_X1 U2615 ( .A(n2240), .ZN(n2305) );
  NOR2_X1 U2616 ( .A1(n2356), .A2(n1873), .ZN(n1958) );
  INV_X1 U2617 ( .A(n1142), .ZN(n2159) );
  NAND2_X1 U2618 ( .A1(mul_operand_b_q[7]), .A2(n2189), .ZN(n2389) );
  AND2_X1 U2619 ( .A1(n2281), .A2(n2282), .ZN(n2392) );
  NOR2_X1 U2620 ( .A1(n2189), .A2(n2191), .ZN(n2390) );
  NAND2_X1 U2621 ( .A1(n2281), .A2(n2390), .ZN(n2391) );
  INV_X1 U2622 ( .A(n2189), .ZN(n2386) );
  INV_X1 U2623 ( .A(mul_operand_b_q[7]), .ZN(n2387) );
  NAND2_X1 U2624 ( .A1(n2386), .A2(n2387), .ZN(n2388) );
  NAND2_X1 U2625 ( .A1(mul_operand_b_q[11]), .A2(mul_operand_b_q[10]), .ZN(
        n2319) );
  AND2_X1 U2626 ( .A1(n2233), .A2(n2244), .ZN(n2322) );
  NOR2_X1 U2627 ( .A1(n2187), .A2(mul_operand_b_q[10]), .ZN(n2320) );
  NAND2_X1 U2628 ( .A1(n2233), .A2(n2320), .ZN(n2321) );
  INV_X1 U2629 ( .A(mul_operand_b_q[10]), .ZN(n2316) );
  INV_X1 U2630 ( .A(mul_operand_b_q[11]), .ZN(n2317) );
  NAND2_X1 U2631 ( .A1(n2316), .A2(n2317), .ZN(n2318) );
  NAND2_X1 U2632 ( .A1(n2321), .A2(n2318), .ZN(n2323) );
  NAND2_X1 U2633 ( .A1(n2323), .A2(n2319), .ZN(n2324) );
  NOR2_X1 U2634 ( .A1(mul_operand_b_q[18]), .A2(mul_operand_b_q[19]), .ZN(
        n2364) );
  AOI21_X1 U2635 ( .B1(n2365), .B2(n2364), .A(n2369), .ZN(n2370) );
  NOR2_X1 U2636 ( .A1(n2364), .A2(n2366), .ZN(n2367) );
  OAI21_X1 U2637 ( .B1(n2365), .B2(n2366), .A(n2414), .ZN(n2368) );
  AOI21_X1 U2638 ( .B1(n2370), .B2(n2429), .A(n2368), .ZN(n2372) );
  INV_X1 U2639 ( .A(n1252), .ZN(n2155) );
  OR2_X1 U2640 ( .A1(n1249), .A2(n2155), .ZN(n2417) );
  INV_X1 U2641 ( .A(mult_x_6_n338), .ZN(n2169) );
  INV_X1 U2642 ( .A(n1147), .ZN(n2157) );
  OR2_X1 U2643 ( .A1(n1144), .A2(n2157), .ZN(n2416) );
  INV_X1 U2644 ( .A(mult_x_6_n350), .ZN(n2163) );
  INV_X1 U2645 ( .A(n1462), .ZN(n2151) );
  OR2_X1 U2646 ( .A1(n1459), .A2(n2151), .ZN(n2419) );
  INV_X1 U2647 ( .A(n1357), .ZN(n2153) );
  OR2_X1 U2648 ( .A1(n1354), .A2(n2153), .ZN(n2418) );
  INV_X1 U2649 ( .A(mult_x_6_n369), .ZN(n2168) );
  BUF_X1 U2650 ( .A(n1246), .Z(n2197) );
  INV_X1 U2651 ( .A(mult_x_6_n393), .ZN(n2162) );
  INV_X1 U2652 ( .A(n1670), .ZN(n2147) );
  OR2_X1 U2653 ( .A1(n1667), .A2(n2147), .ZN(n2426) );
  BUF_X1 U2654 ( .A(mul_operand_b_q[16]), .Z(n2184) );
  INV_X1 U2655 ( .A(n1567), .ZN(n2149) );
  OR2_X1 U2656 ( .A1(n1564), .A2(n2149), .ZN(n2425) );
  BUF_X1 U2657 ( .A(n1351), .Z(n2199) );
  INV_X1 U2658 ( .A(mult_x_6_n424), .ZN(n2167) );
  INV_X1 U2659 ( .A(mult_x_6_n460), .ZN(n2161) );
  XNOR2_X1 U2660 ( .A(mul_operand_a_q[5]), .B(mul_operand_a_q[6]), .ZN(n1873)
         );
  INV_X1 U2661 ( .A(n18701), .ZN(n2342) );
  NAND2_X1 U2662 ( .A1(n1873), .A2(n2342), .ZN(n2215) );
  BUF_X1 U2663 ( .A(mul_operand_b_q[9]), .Z(n2186) );
  INV_X1 U2664 ( .A(n1769), .ZN(n2406) );
  NAND2_X1 U2665 ( .A1(n1772), .A2(n2406), .ZN(n2210) );
  INV_X1 U2666 ( .A(n2418), .ZN(n2200) );
  INV_X1 U2667 ( .A(mult_x_6_n503), .ZN(n2166) );
  INV_X1 U2668 ( .A(mult_x_6_n551), .ZN(n2160) );
  BUF_X1 U2669 ( .A(n1560), .Z(n2201) );
  INV_X1 U2670 ( .A(mult_x_6_n664), .ZN(n2164) );
  INV_X1 U2671 ( .A(n2049), .ZN(n2143) );
  INV_X1 U2672 ( .A(n2144), .ZN(n2329) );
  NAND3_X1 U2673 ( .A1(n2329), .A2(n2143), .A3(n2427), .ZN(n1961) );
  BUF_X1 U2674 ( .A(mul_operand_b_q[5]), .Z(n2190) );
  INV_X1 U2675 ( .A(mult_x_6_n606), .ZN(n2165) );
  BUF_X1 U2676 ( .A(mul_operand_b_q[6]), .Z(n2188) );
  BUF_X1 U2677 ( .A(mul_operand_b_q[1]), .Z(n2286) );
  BUF_X1 U2678 ( .A(n1768), .Z(n2208) );
  BUF_X1 U2679 ( .A(n1869), .Z(n2212) );
  INV_X1 U2680 ( .A(n2210), .ZN(n2211) );
  INV_X1 U2681 ( .A(n2426), .ZN(n2206) );
  INV_X1 U2682 ( .A(n1874), .ZN(n2356) );
  INV_X1 U2683 ( .A(n1875), .ZN(n2145) );
  NAND2_X1 U2684 ( .A1(mult_x_6_n817), .A2(mult_x_6_n1395), .ZN(n2397) );
  NAND2_X1 U2685 ( .A1(mult_x_6_n731), .A2(mult_x_6_n1390), .ZN(n2384) );
  INV_X1 U2686 ( .A(mult_x_6_n1386), .ZN(n2377) );
  XNOR2_X1 U2687 ( .A(mult_x_6_n651), .B(n2377), .ZN(n2378) );
  XNOR2_X1 U2688 ( .A(n2378), .B(n2379), .ZN(mult_x_6_n649) );
  BUF_X1 U2689 ( .A(n2048), .Z(n2222) );
  XNOR2_X1 U2690 ( .A(mult_x_6_n731), .B(mult_x_6_n1390), .ZN(n2383) );
  XNOR2_X1 U2691 ( .A(mult_x_6_n817), .B(mult_x_6_n1395), .ZN(n2396) );
  NAND2_X1 U2692 ( .A1(mult_x_6_n845), .A2(mult_x_6_n1429), .ZN(n2327) );
  XNOR2_X1 U2693 ( .A(n2034), .B(n1026), .ZN(n2359) );
  NAND2_X1 U2694 ( .A1(mult_x_6_n1443), .A2(mult_x_6_n981), .ZN(n2403) );
  XNOR2_X1 U2695 ( .A(mult_x_6_n941), .B(mult_x_6_n1405), .ZN(n2400) );
  NAND2_X1 U2696 ( .A1(n2359), .A2(mult_x_6_n947), .ZN(n2355) );
  XNOR2_X1 U2697 ( .A(mult_x_6_n671), .B(mult_x_6_n1387), .ZN(n2363) );
  NOR2_X1 U2698 ( .A1(n1014), .A2(mul_operand_a_q[0]), .ZN(n2141) );
  NOR2_X1 U2699 ( .A1(n2399), .A2(n2405), .ZN(n2120) );
  XNOR2_X1 U2700 ( .A(mult_x_6_n799), .B(mult_x_6_n1426), .ZN(n2349) );
  XNOR2_X1 U2701 ( .A(mult_x_6_n845), .B(mult_x_6_n1429), .ZN(n2326) );
  XNOR2_X1 U2702 ( .A(mult_x_6_n859), .B(mult_x_6_n1430), .ZN(n2330) );
  NAND2_X1 U2703 ( .A1(n2360), .A2(n2355), .ZN(n2357) );
  XNOR2_X1 U2704 ( .A(mult_x_6_n939), .B(mult_x_6_n1437), .ZN(n2358) );
  XNOR2_X1 U2705 ( .A(mult_x_6_n1443), .B(mult_x_6_n981), .ZN(n2402) );
  OR2_X1 U2706 ( .A1(mult_x_6_n979), .A2(mult_x_6_n1475), .ZN(n2398) );
  XNOR2_X1 U2707 ( .A(mult_x_6_n669), .B(mult_x_6_n1419), .ZN(n2344) );
  NOR2_X1 U2708 ( .A1(mult_x_6_n609), .A2(mult_x_6_n627), .ZN(n2331) );
  NOR2_X1 U2709 ( .A1(mult_x_6_n554), .A2(mult_x_6_n570), .ZN(n2334) );
  NOR2_X1 U2710 ( .A1(mult_x_6_n535), .A2(mult_x_6_n521), .ZN(n2338) );
  NOR2_X1 U2711 ( .A1(mult_x_6_n505), .A2(mult_x_6_n490), .ZN(n2343) );
  NOR2_X1 U2712 ( .A1(mult_x_6_n462), .A2(mult_x_6_n449), .ZN(n2288) );
  NOR2_X1 U2713 ( .A1(n2289), .A2(n2430), .ZN(n2293) );
  INV_X1 U2714 ( .A(mult_x_6_n438), .ZN(n2294) );
  NOR2_X1 U2715 ( .A1(n2293), .A2(n2294), .ZN(n2295) );
  INV_X1 U2716 ( .A(mult_x_6_n448), .ZN(n2290) );
  NOR2_X1 U2717 ( .A1(n2288), .A2(n2290), .ZN(n2291) );
  NOR2_X1 U2718 ( .A1(n2295), .A2(n2291), .ZN(n2297) );
  AOI21_X1 U2719 ( .B1(n2295), .B2(n2430), .A(n2292), .ZN(n2298) );
  NOR2_X1 U2720 ( .A1(mult_x_6_n395), .A2(mult_x_6_n386), .ZN(n2336) );
  NOR2_X1 U2721 ( .A1(mult_x_6_n371), .A2(mult_x_6_n364), .ZN(n2333) );
  NOR2_X1 U2722 ( .A1(mult_x_6_n353), .A2(mult_x_6_n357), .ZN(n2337) );
  NOR2_X1 U2723 ( .A1(mult_x_6_n346), .A2(mult_x_6_n344), .ZN(n2299) );
  INV_X1 U2724 ( .A(n2299), .ZN(n2300) );
  OAI21_X1 U2725 ( .B1(n2254), .B2(n2300), .A(mult_x_6_n343), .ZN(n2301) );
  INV_X1 U2726 ( .A(n2301), .ZN(n2302) );
  INV_X1 U2727 ( .A(mult_x_6_n333), .ZN(n2304) );
  INV_X1 U2728 ( .A(mult_x_6_n334), .ZN(n2306) );
  AOI21_X1 U2729 ( .B1(n2310), .B2(n2240), .A(n2306), .ZN(n2307) );
  NOR2_X1 U2730 ( .A1(mult_x_6_n336), .A2(mult_x_6_n335), .ZN(n2310) );
  NAND2_X1 U2731 ( .A1(n2240), .A2(n2310), .ZN(n2312) );
  AOI22_X1 U2732 ( .A1(n2242), .A2(n2312), .B1(n2309), .B2(n2240), .ZN(n2313)
         );
  INV_X1 U2733 ( .A(n2310), .ZN(n2311) );
  AOI21_X1 U2734 ( .B1(mult_x_6_n286), .B2(n2289), .A(n2430), .ZN(n2296) );
  INV_X1 U2735 ( .A(n2296), .ZN(mult_x_6_n285) );
  BUF_X2 U2736 ( .A(mul_operand_b_q[30]), .Z(n2180) );
  BUF_X2 U2737 ( .A(mul_operand_a_q[20]), .Z(n2170) );
  BUF_X2 U2738 ( .A(mul_operand_a_q[14]), .Z(n2172) );
  BUF_X2 U2739 ( .A(mul_operand_a_q[17]), .Z(n2171) );
  BUF_X2 U2740 ( .A(mul_operand_a_q[11]), .Z(n2173) );
  BUF_X1 U2741 ( .A(mul_operand_b_q[32]), .Z(n2177) );
  BUF_X1 U2742 ( .A(n1958), .Z(n2213) );
  BUF_X1 U2743 ( .A(mul_operand_b_q[28]), .Z(n2181) );
  BUF_X1 U2744 ( .A(mul_operand_b_q[26]), .Z(n2182) );
  AND2_X1 U2745 ( .A1(mul_operand_b_q[19]), .A2(mul_operand_b_q[18]), .ZN(
        n2429) );
  BUF_X1 U2746 ( .A(mul_operand_b_q[24]), .Z(n2183) );
  BUF_X1 U2747 ( .A(mul_operand_b_q[16]), .Z(n2185) );
  NAND2_X1 U2748 ( .A1(mult_x_6_n1064), .A2(mul_operand_b_q[8]), .ZN(n2253) );
  NAND2_X1 U2749 ( .A1(mult_x_6_n1064), .A2(mul_operand_b_q[7]), .ZN(n2252) );
  NAND2_X1 U2750 ( .A1(n2250), .A2(mul_operand_b_q[23]), .ZN(n2236) );
  AND2_X1 U2751 ( .A1(mult_x_6_n449), .A2(mult_x_6_n462), .ZN(n2430) );
  AND2_X1 U2752 ( .A1(n2196), .A2(mul_operand_a_q[0]), .ZN(n2431) );
  NAND3_X1 U2753 ( .A1(n2434), .A2(n2433), .A3(n2432), .ZN(mult_x_6_n327) );
  NAND2_X1 U2754 ( .A1(mult_x_6_n1480), .A2(mult_x_6_n995), .ZN(n2432) );
  NAND2_X1 U2755 ( .A1(mult_x_6_n328), .A2(mult_x_6_n995), .ZN(n2433) );
  NAND2_X1 U2756 ( .A1(mult_x_6_n1480), .A2(mult_x_6_n328), .ZN(n2434) );
  XOR2_X1 U2757 ( .A(mult_x_6_n328), .B(n2435), .Z(mult_result_w[3]) );
  XOR2_X1 U2758 ( .A(mult_x_6_n1480), .B(mult_x_6_n995), .Z(n2435) );
  NAND2_X1 U2759 ( .A1(mult_x_6_n843), .A2(mult_x_6_n1461), .ZN(n2436) );
  XOR2_X1 U2760 ( .A(mult_x_6_n309), .B(n2437), .Z(mult_result_w[22]) );
  XOR2_X1 U2761 ( .A(mult_x_6_n843), .B(mult_x_6_n1461), .Z(n2437) );
  XOR2_X1 U2762 ( .A(n1027), .B(n2438), .Z(mult_result_w[43]) );
  XOR2_X1 U2763 ( .A(mult_x_6_n489), .B(mult_x_6_n476), .Z(n2438) );
  BUF_X2 U2764 ( .A(n2048), .Z(n2223) );
  XOR2_X1 U2765 ( .A(n2439), .B(n1013), .Z(mult_x_6_n1478) );
  XOR2_X1 U2766 ( .A(mult_x_6_n966), .B(n2440), .Z(mult_x_6_n961) );
  XOR2_X1 U2767 ( .A(mult_x_6_n1440), .B(mult_x_6_n963), .Z(n2440) );
  XOR2_X1 U2768 ( .A(mult_x_6_n1447), .B(mult_x_6_n994), .Z(mult_x_6_n993) );
  XNOR2_X1 U2769 ( .A(n1009), .B(n2194), .ZN(n2441) );
  NOR2_X2 U2770 ( .A1(n2973), .A2(n2473), .ZN(n2801) );
  BUF_X1 U2771 ( .A(n2742), .Z(n2568) );
  INV_X1 U2772 ( .A(n2969), .ZN(n2803) );
  BUF_X1 U2773 ( .A(n2744), .Z(n2569) );
  BUF_X1 U2774 ( .A(n2745), .Z(n2570) );
  OR2_X1 U2775 ( .A1(n2804), .A2(n2817), .ZN(n2499) );
  BUF_X1 U2776 ( .A(n2882), .Z(n2576) );
  BUF_X1 U2777 ( .A(n2881), .Z(n2575) );
  BUF_X1 U2778 ( .A(n2967), .Z(n2577) );
  NAND2_X1 U2779 ( .A1(n2966), .A2(n2574), .ZN(n2742) );
  NAND2_X1 U2780 ( .A1(n2802), .A2(n2803), .ZN(n2971) );
  AOI21_X1 U2781 ( .B1(n2818), .B2(n2822), .A(n2821), .ZN(n2969) );
  NOR2_X1 U2782 ( .A1(n2574), .A2(n2968), .ZN(n2741) );
  NOR2_X1 U2783 ( .A1(n2819), .A2(n2803), .ZN(n2881) );
  INV_X1 U2784 ( .A(n2971), .ZN(n2968) );
  BUF_X1 U2785 ( .A(n2800), .Z(n2571) );
  BUF_X1 U2786 ( .A(n2994), .Z(n2579) );
  BUF_X1 U2787 ( .A(n2993), .Z(n2578) );
  INV_X1 U2788 ( .A(rst_i), .ZN(n2802) );
  INV_X1 U2789 ( .A(operand_rb_i[31]), .ZN(n2820) );
  BUF_X2 U2790 ( .A(n2801), .Z(n2574) );
  NAND2_X1 U2791 ( .A1(n2972), .A2(n2802), .ZN(n2973) );
  NOR2_X1 U2792 ( .A1(n2975), .A2(n104), .ZN(n2800) );
  INV_X2 U2793 ( .A(n2486), .ZN(n2580) );
  INV_X2 U2794 ( .A(n2487), .ZN(n2581) );
  NOR3_X1 U2795 ( .A1(mulhi_sel_q), .A2(n2470), .A3(n2973), .ZN(n2994) );
  NOR3_X1 U2796 ( .A1(n2973), .A2(n2470), .A3(n2526), .ZN(n2993) );
  NAND2_X1 U2797 ( .A1(n2803), .A2(n2573), .ZN(n578) );
  OAI21_X1 U2798 ( .B1(n2971), .B2(n2483), .A(n2970), .ZN(n449) );
  AOI21_X1 U2799 ( .B1(n406), .B2(divisor_q[16]), .A(n2658), .ZN(n305) );
  INV_X1 U2800 ( .A(n2657), .ZN(n2658) );
  AOI21_X1 U2801 ( .B1(n406), .B2(divisor_q[0]), .A(n2706), .ZN(n321) );
  INV_X1 U2802 ( .A(n2705), .ZN(n2706) );
  AOI21_X1 U2803 ( .B1(n406), .B2(divisor_q[15]), .A(n2661), .ZN(n306) );
  INV_X1 U2804 ( .A(n2660), .ZN(n2661) );
  AOI21_X1 U2805 ( .B1(n406), .B2(divisor_q[11]), .A(n2673), .ZN(n310) );
  INV_X1 U2806 ( .A(n2672), .ZN(n2673) );
  AOI21_X1 U2807 ( .B1(n406), .B2(divisor_q[22]), .A(n2640), .ZN(n299) );
  INV_X1 U2808 ( .A(n2639), .ZN(n2640) );
  AOI21_X1 U2809 ( .B1(n406), .B2(divisor_q[18]), .A(n2652), .ZN(n303) );
  INV_X1 U2810 ( .A(n2651), .ZN(n2652) );
  AOI21_X1 U2811 ( .B1(n406), .B2(divisor_q[17]), .A(n2655), .ZN(n304) );
  INV_X1 U2812 ( .A(n2654), .ZN(n2655) );
  OAI22_X1 U2813 ( .A1(n2742), .A2(n6400), .B1(n96), .B2(n2741), .ZN(n473) );
  OAI22_X1 U2814 ( .A1(n2742), .A2(n2519), .B1(n99), .B2(n2741), .ZN(n476) );
  OAI22_X1 U2815 ( .A1(n2742), .A2(n2518), .B1(n97), .B2(n2741), .ZN(n474) );
  OAI22_X1 U2816 ( .A1(n2742), .A2(n2465), .B1(n95), .B2(n2741), .ZN(n472) );
  AOI21_X1 U2817 ( .B1(n406), .B2(divisor_q[27]), .A(n2625), .ZN(n294) );
  INV_X1 U2818 ( .A(n2624), .ZN(n2625) );
  AOI21_X1 U2819 ( .B1(n406), .B2(divisor_q[1]), .A(n2703), .ZN(n320) );
  INV_X1 U2820 ( .A(n2702), .ZN(n2703) );
  AOI21_X1 U2821 ( .B1(n406), .B2(divisor_q[23]), .A(n2637), .ZN(n298) );
  INV_X1 U2822 ( .A(n2636), .ZN(n2637) );
  AOI21_X1 U2823 ( .B1(n406), .B2(divisor_q[25]), .A(n2631), .ZN(n296) );
  INV_X1 U2824 ( .A(n2630), .ZN(n2631) );
  AOI21_X1 U2825 ( .B1(n406), .B2(divisor_q[24]), .A(n2634), .ZN(n297) );
  INV_X1 U2826 ( .A(n2633), .ZN(n2634) );
  AOI21_X1 U2827 ( .B1(n406), .B2(divisor_q[28]), .A(n2622), .ZN(n293) );
  INV_X1 U2828 ( .A(n2621), .ZN(n2622) );
  AOI21_X1 U2829 ( .B1(n406), .B2(divisor_q[21]), .A(n2643), .ZN(n300) );
  INV_X1 U2830 ( .A(n2642), .ZN(n2643) );
  AOI21_X1 U2831 ( .B1(n406), .B2(divisor_q[26]), .A(n2628), .ZN(n295) );
  INV_X1 U2832 ( .A(n2627), .ZN(n2628) );
  AOI21_X1 U2833 ( .B1(n406), .B2(divisor_q[29]), .A(n2619), .ZN(n292) );
  INV_X1 U2834 ( .A(n2618), .ZN(n2619) );
  AOI21_X1 U2835 ( .B1(n406), .B2(divisor_q[13]), .A(n2667), .ZN(n308) );
  INV_X1 U2836 ( .A(n2666), .ZN(n2667) );
  AOI21_X1 U2837 ( .B1(n406), .B2(divisor_q[20]), .A(n2646), .ZN(n301) );
  INV_X1 U2838 ( .A(n2645), .ZN(n2646) );
  AOI21_X1 U2839 ( .B1(n406), .B2(divisor_q[19]), .A(n2649), .ZN(n302) );
  INV_X1 U2840 ( .A(n2648), .ZN(n2649) );
  AOI21_X1 U2841 ( .B1(n406), .B2(divisor_q[14]), .A(n2664), .ZN(n307) );
  INV_X1 U2842 ( .A(n2663), .ZN(n2664) );
  AOI21_X1 U2843 ( .B1(n406), .B2(divisor_q[2]), .A(n2700), .ZN(n319) );
  INV_X1 U2844 ( .A(n2699), .ZN(n2700) );
  AOI21_X1 U2845 ( .B1(n406), .B2(divisor_q[9]), .A(n2679), .ZN(n312) );
  INV_X1 U2846 ( .A(n2678), .ZN(n2679) );
  AOI21_X1 U2847 ( .B1(n406), .B2(divisor_q[3]), .A(n2697), .ZN(n318) );
  INV_X1 U2848 ( .A(n2696), .ZN(n2697) );
  AOI21_X1 U2849 ( .B1(n406), .B2(divisor_q[12]), .A(n2670), .ZN(n309) );
  INV_X1 U2850 ( .A(n2669), .ZN(n2670) );
  AOI21_X1 U2851 ( .B1(n406), .B2(divisor_q[5]), .A(n2691), .ZN(n316) );
  INV_X1 U2852 ( .A(n2690), .ZN(n2691) );
  AOI21_X1 U2853 ( .B1(n406), .B2(divisor_q[6]), .A(n2688), .ZN(n315) );
  INV_X1 U2854 ( .A(n2687), .ZN(n2688) );
  AOI21_X1 U2855 ( .B1(n406), .B2(divisor_q[7]), .A(n2685), .ZN(n314) );
  INV_X1 U2856 ( .A(n2684), .ZN(n2685) );
  AOI21_X1 U2857 ( .B1(n406), .B2(divisor_q[8]), .A(n2682), .ZN(n313) );
  INV_X1 U2858 ( .A(n2681), .ZN(n2682) );
  AOI21_X1 U2859 ( .B1(n406), .B2(divisor_q[4]), .A(n2694), .ZN(n317) );
  INV_X1 U2860 ( .A(n2693), .ZN(n2694) );
  AOI21_X1 U2861 ( .B1(n406), .B2(divisor_q[10]), .A(n2676), .ZN(n311) );
  INV_X1 U2862 ( .A(n2675), .ZN(n2676) );
  OAI21_X1 U2863 ( .B1(n2803), .B2(n2535), .A(n2614), .ZN(n544) );
  AOI22_X1 U2864 ( .A1(n406), .A2(divisor_q[31]), .B1(n2574), .B2(
        divisor_q[32]), .ZN(n2614) );
  AOI21_X1 U2865 ( .B1(divisor_q[30]), .B2(n406), .A(n2616), .ZN(n290) );
  INV_X1 U2866 ( .A(n2615), .ZN(n2616) );
  OAI22_X1 U2867 ( .A1(n2742), .A2(n2458), .B1(n98), .B2(n6101), .ZN(n475) );
  OAI22_X1 U2868 ( .A1(n2742), .A2(n2446), .B1(n101), .B2(n6101), .ZN(n478) );
  OAI22_X1 U2869 ( .A1(n2742), .A2(n2516), .B1(n8100), .B2(n6101), .ZN(n458)
         );
  OAI22_X1 U2870 ( .A1(n2742), .A2(n2466), .B1(n8500), .B2(n6101), .ZN(n462)
         );
  OAI22_X1 U2871 ( .A1(n2742), .A2(n2521), .B1(n8400), .B2(n6101), .ZN(n461)
         );
  OAI22_X1 U2872 ( .A1(n2742), .A2(n2523), .B1(n102), .B2(n6101), .ZN(n479) );
  OAI22_X1 U2873 ( .A1(n2742), .A2(n2460), .B1(n8000), .B2(n6101), .ZN(n457)
         );
  OAI22_X1 U2874 ( .A1(n2742), .A2(n2464), .B1(n100), .B2(n6101), .ZN(n477) );
  OAI22_X1 U2875 ( .A1(n2742), .A2(n2467), .B1(n8200), .B2(n6101), .ZN(n459)
         );
  OAI22_X1 U2876 ( .A1(n2742), .A2(n2445), .B1(n8300), .B2(n6101), .ZN(n460)
         );
  OAI22_X1 U2877 ( .A1(n2742), .A2(n2513), .B1(n7900), .B2(n6101), .ZN(n456)
         );
  OAI22_X1 U2878 ( .A1(n2568), .A2(n2512), .B1(n8600), .B2(n6101), .ZN(n463)
         );
  OAI22_X1 U2879 ( .A1(n2568), .A2(n2515), .B1(n7400), .B2(n6101), .ZN(n451)
         );
  OAI22_X1 U2880 ( .A1(n2568), .A2(n2461), .B1(n7300), .B2(n6101), .ZN(n450)
         );
  OAI22_X1 U2881 ( .A1(n2568), .A2(n2469), .B1(n90), .B2(n6101), .ZN(n467) );
  OAI22_X1 U2882 ( .A1(n2568), .A2(n2517), .B1(n8900), .B2(n6101), .ZN(n466)
         );
  OAI22_X1 U2883 ( .A1(n2568), .A2(n2443), .B1(n8800), .B2(n6101), .ZN(n465)
         );
  OAI22_X1 U2884 ( .A1(n2568), .A2(n2459), .B1(n87), .B2(n6101), .ZN(n464) );
  OAI22_X1 U2885 ( .A1(n2568), .A2(n2444), .B1(n7600), .B2(n6101), .ZN(n453)
         );
  OAI22_X1 U2886 ( .A1(n2568), .A2(n2468), .B1(n7800), .B2(n6101), .ZN(n455)
         );
  OAI22_X1 U2887 ( .A1(n2568), .A2(n2522), .B1(n7700), .B2(n6101), .ZN(n454)
         );
  OAI22_X1 U2888 ( .A1(n2568), .A2(n7100), .B1(n103), .B2(n6101), .ZN(n480) );
  OAI22_X1 U2889 ( .A1(n2568), .A2(n2463), .B1(n7500), .B2(n6101), .ZN(n452)
         );
  OAI22_X1 U2890 ( .A1(n2568), .A2(n2514), .B1(n91), .B2(n6101), .ZN(n468) );
  OAI22_X1 U2891 ( .A1(n2568), .A2(n2462), .B1(n92), .B2(n6101), .ZN(n469) );
  OAI22_X1 U2892 ( .A1(n2568), .A2(n2511), .B1(n7200), .B2(n6101), .ZN(n481)
         );
  OAI22_X1 U2893 ( .A1(n2568), .A2(n2442), .B1(n93), .B2(n6101), .ZN(n470) );
  OAI22_X1 U2894 ( .A1(n2568), .A2(n2520), .B1(n94), .B2(n6101), .ZN(n471) );
  INV_X1 U2895 ( .A(n2611), .ZN(n510) );
  INV_X1 U2896 ( .A(n2612), .ZN(n511) );
  INV_X1 U2897 ( .A(n2613), .ZN(n512) );
  AOI222_X1 U2898 ( .A1(n2710), .A2(C21_DATA3_0), .B1(n2709), .B2(
        operand_ra_i[0]), .C1(dividend_q[0]), .C2(n2577), .ZN(n2613) );
  INV_X1 U2899 ( .A(n2610), .ZN(n509) );
  AOI222_X1 U2900 ( .A1(n2710), .A2(C21_DATA3_3), .B1(n2709), .B2(
        operand_ra_i[3]), .C1(dividend_q[3]), .C2(n2577), .ZN(n2610) );
  INV_X1 U2901 ( .A(n2608), .ZN(n507) );
  AOI222_X1 U2902 ( .A1(n2710), .A2(C21_DATA3_5), .B1(n2709), .B2(
        operand_ra_i[5]), .C1(dividend_q[5]), .C2(n2577), .ZN(n2608) );
  INV_X1 U2903 ( .A(n2605), .ZN(n504) );
  AOI222_X1 U2904 ( .A1(n2710), .A2(C21_DATA3_8), .B1(n2709), .B2(
        operand_ra_i[8]), .C1(dividend_q[8]), .C2(n2577), .ZN(n2605) );
  INV_X1 U2905 ( .A(n2609), .ZN(n508) );
  AOI222_X1 U2906 ( .A1(n2710), .A2(C21_DATA3_4), .B1(n2709), .B2(
        operand_ra_i[4]), .C1(dividend_q[4]), .C2(n2577), .ZN(n2609) );
  INV_X1 U2907 ( .A(n2607), .ZN(n506) );
  AOI222_X1 U2908 ( .A1(n2710), .A2(C21_DATA3_6), .B1(n2709), .B2(
        operand_ra_i[6]), .C1(dividend_q[6]), .C2(n2577), .ZN(n2607) );
  INV_X1 U2909 ( .A(n2606), .ZN(n505) );
  AOI222_X1 U2910 ( .A1(n2710), .A2(C21_DATA3_7), .B1(n2709), .B2(
        operand_ra_i[7]), .C1(dividend_q[7]), .C2(n2967), .ZN(n2606) );
  INV_X1 U2911 ( .A(n2604), .ZN(n503) );
  AOI222_X1 U2912 ( .A1(n2710), .A2(C21_DATA3_9), .B1(n2709), .B2(
        operand_ra_i[9]), .C1(dividend_q[9]), .C2(n2577), .ZN(n2604) );
  INV_X1 U2913 ( .A(n2603), .ZN(n502) );
  AOI222_X1 U2914 ( .A1(n2710), .A2(C21_DATA3_10), .B1(n2709), .B2(
        operand_ra_i[10]), .C1(dividend_q[10]), .C2(n2577), .ZN(n2603) );
  INV_X1 U2915 ( .A(n2602), .ZN(n501) );
  AOI222_X1 U2916 ( .A1(n2710), .A2(C21_DATA3_11), .B1(n2709), .B2(
        operand_ra_i[11]), .C1(dividend_q[11]), .C2(n2967), .ZN(n2602) );
  INV_X1 U2917 ( .A(operand_rb_i[30]), .ZN(n2565) );
  INV_X1 U2918 ( .A(operand_rb_i[29]), .ZN(n2564) );
  INV_X1 U2919 ( .A(operand_rb_i[28]), .ZN(n2563) );
  INV_X1 U2920 ( .A(operand_rb_i[27]), .ZN(n2562) );
  INV_X1 U2921 ( .A(operand_rb_i[26]), .ZN(n2561) );
  INV_X1 U2922 ( .A(operand_rb_i[25]), .ZN(n2560) );
  INV_X1 U2923 ( .A(operand_rb_i[24]), .ZN(n2559) );
  INV_X1 U2924 ( .A(operand_rb_i[23]), .ZN(n2558) );
  INV_X1 U2925 ( .A(operand_rb_i[22]), .ZN(n2557) );
  INV_X1 U2926 ( .A(operand_rb_i[21]), .ZN(n2556) );
  INV_X1 U2927 ( .A(operand_rb_i[20]), .ZN(n2555) );
  INV_X1 U2928 ( .A(operand_rb_i[19]), .ZN(n2554) );
  INV_X1 U2929 ( .A(operand_rb_i[18]), .ZN(n2553) );
  INV_X1 U2930 ( .A(operand_rb_i[17]), .ZN(n2552) );
  INV_X1 U2931 ( .A(operand_rb_i[16]), .ZN(n2551) );
  INV_X1 U2932 ( .A(operand_rb_i[15]), .ZN(n2550) );
  INV_X1 U2933 ( .A(operand_rb_i[14]), .ZN(n2549) );
  INV_X1 U2934 ( .A(operand_rb_i[13]), .ZN(n2548) );
  INV_X1 U2935 ( .A(operand_rb_i[12]), .ZN(n2547) );
  INV_X1 U2936 ( .A(operand_rb_i[11]), .ZN(n2546) );
  INV_X1 U2937 ( .A(operand_rb_i[10]), .ZN(n2545) );
  INV_X1 U2938 ( .A(operand_rb_i[9]), .ZN(n2544) );
  INV_X1 U2939 ( .A(operand_rb_i[8]), .ZN(n2543) );
  INV_X1 U2940 ( .A(operand_rb_i[7]), .ZN(n2542) );
  INV_X1 U2941 ( .A(operand_rb_i[6]), .ZN(n2541) );
  INV_X1 U2942 ( .A(operand_rb_i[5]), .ZN(n2540) );
  INV_X1 U2943 ( .A(operand_rb_i[4]), .ZN(n2539) );
  INV_X1 U2944 ( .A(operand_rb_i[3]), .ZN(n2538) );
  INV_X1 U2945 ( .A(operand_rb_i[2]), .ZN(n2537) );
  INV_X1 U2946 ( .A(n2601), .ZN(n500) );
  AOI222_X1 U2947 ( .A1(n2710), .A2(C21_DATA3_12), .B1(n2709), .B2(
        operand_ra_i[12]), .C1(dividend_q[12]), .C2(n2577), .ZN(n2601) );
  INV_X1 U2948 ( .A(n2600), .ZN(n499) );
  AOI222_X1 U2949 ( .A1(n2710), .A2(C21_DATA3_13), .B1(n2709), .B2(
        operand_ra_i[13]), .C1(dividend_q[13]), .C2(n2577), .ZN(n2600) );
  INV_X1 U2950 ( .A(n2599), .ZN(n498) );
  AOI222_X1 U2951 ( .A1(n2710), .A2(C21_DATA3_14), .B1(n2709), .B2(
        operand_ra_i[14]), .C1(dividend_q[14]), .C2(n2967), .ZN(n2599) );
  INV_X1 U2952 ( .A(n2598), .ZN(n497) );
  AOI222_X1 U2953 ( .A1(n2710), .A2(C21_DATA3_15), .B1(n2709), .B2(
        operand_ra_i[15]), .C1(dividend_q[15]), .C2(n2577), .ZN(n2598) );
  INV_X1 U2954 ( .A(n2597), .ZN(n496) );
  AOI222_X1 U2955 ( .A1(n2710), .A2(C21_DATA3_16), .B1(n2709), .B2(
        operand_ra_i[16]), .C1(dividend_q[16]), .C2(n2967), .ZN(n2597) );
  INV_X1 U2956 ( .A(n2596), .ZN(n495) );
  AOI222_X1 U2957 ( .A1(n2710), .A2(C21_DATA3_17), .B1(n2709), .B2(
        operand_ra_i[17]), .C1(dividend_q[17]), .C2(n2577), .ZN(n2596) );
  INV_X1 U2958 ( .A(n2595), .ZN(n494) );
  AOI222_X1 U2959 ( .A1(n2710), .A2(C21_DATA3_18), .B1(n2709), .B2(
        operand_ra_i[18]), .C1(dividend_q[18]), .C2(n2577), .ZN(n2595) );
  INV_X1 U2960 ( .A(n2594), .ZN(n493) );
  AOI222_X1 U2961 ( .A1(n2710), .A2(C21_DATA3_19), .B1(n2709), .B2(
        operand_ra_i[19]), .C1(dividend_q[19]), .C2(n2967), .ZN(n2594) );
  INV_X1 U2962 ( .A(n2593), .ZN(n492) );
  AOI222_X1 U2963 ( .A1(n2710), .A2(C21_DATA3_20), .B1(n2709), .B2(
        operand_ra_i[20]), .C1(dividend_q[20]), .C2(n2967), .ZN(n2593) );
  NAND2_X1 U2964 ( .A1(n2992), .A2(n2750), .ZN(n420) );
  AOI21_X1 U2965 ( .B1(n2800), .B2(C22_DATA3_3), .A(n2749), .ZN(n2750) );
  OAI21_X1 U2966 ( .B1(n2799), .B2(n100), .A(n2748), .ZN(n2749) );
  AOI22_X1 U2967 ( .A1(n2581), .A2(dividend_q[3]), .B1(result_o[3]), .B2(n2580), .ZN(n2748) );
  INV_X1 U2968 ( .A(n2592), .ZN(n491) );
  AOI222_X1 U2969 ( .A1(n2710), .A2(C21_DATA3_21), .B1(n2709), .B2(
        operand_ra_i[21]), .C1(dividend_q[21]), .C2(n2967), .ZN(n2592) );
  NAND2_X1 U2970 ( .A1(n2991), .A2(n2753), .ZN(n421) );
  AOI21_X1 U2971 ( .B1(n2800), .B2(C22_DATA3_4), .A(n2752), .ZN(n2753) );
  OAI21_X1 U2972 ( .B1(n2799), .B2(n99), .A(n2751), .ZN(n2752) );
  AOI22_X1 U2973 ( .A1(result_o[4]), .A2(n2580), .B1(dividend_q[4]), .B2(n2581), .ZN(n2751) );
  INV_X1 U2974 ( .A(n2591), .ZN(n490) );
  AOI222_X1 U2975 ( .A1(n2710), .A2(C21_DATA3_22), .B1(n2709), .B2(
        operand_ra_i[22]), .C1(dividend_q[22]), .C2(n2967), .ZN(n2591) );
  NAND2_X1 U2976 ( .A1(n2990), .A2(n2756), .ZN(n423) );
  AOI21_X1 U2977 ( .B1(C22_DATA3_6), .B2(n2800), .A(n2755), .ZN(n2756) );
  OAI21_X1 U2978 ( .B1(n2799), .B2(n97), .A(n2754), .ZN(n2755) );
  AOI22_X1 U2979 ( .A1(result_o[6]), .A2(n2580), .B1(dividend_q[6]), .B2(n2581), .ZN(n2754) );
  INV_X1 U2980 ( .A(n2590), .ZN(n489) );
  AOI222_X1 U2981 ( .A1(n2710), .A2(C21_DATA3_23), .B1(n2709), .B2(
        operand_ra_i[23]), .C1(dividend_q[23]), .C2(n2967), .ZN(n2590) );
  NAND2_X1 U2982 ( .A1(n2989), .A2(n2759), .ZN(n424) );
  AOI21_X1 U2983 ( .B1(C22_DATA3_7), .B2(n2800), .A(n2758), .ZN(n2759) );
  OAI21_X1 U2984 ( .B1(n2799), .B2(n96), .A(n2757), .ZN(n2758) );
  AOI22_X1 U2985 ( .A1(n2581), .A2(dividend_q[7]), .B1(result_o[7]), .B2(n2580), .ZN(n2757) );
  INV_X1 U2986 ( .A(n2589), .ZN(n488) );
  AOI222_X1 U2987 ( .A1(n2710), .A2(C21_DATA3_24), .B1(n2709), .B2(
        operand_ra_i[24]), .C1(dividend_q[24]), .C2(n2967), .ZN(n2589) );
  INV_X1 U2988 ( .A(n2588), .ZN(n487) );
  AOI222_X1 U2989 ( .A1(n2710), .A2(C21_DATA3_25), .B1(n2709), .B2(
        operand_ra_i[25]), .C1(dividend_q[25]), .C2(n2577), .ZN(n2588) );
  INV_X1 U2990 ( .A(n2587), .ZN(n486) );
  AOI222_X1 U2991 ( .A1(n2710), .A2(C21_DATA3_26), .B1(n2709), .B2(
        operand_ra_i[26]), .C1(dividend_q[26]), .C2(n2967), .ZN(n2587) );
  NAND2_X1 U2992 ( .A1(n2988), .A2(n2762), .ZN(n427) );
  AOI21_X1 U2993 ( .B1(C22_DATA3_10), .B2(n2571), .A(n2761), .ZN(n2762) );
  OAI21_X1 U2994 ( .B1(n2799), .B2(n93), .A(n2760), .ZN(n2761) );
  AOI22_X1 U2995 ( .A1(result_o[10]), .A2(n2580), .B1(dividend_q[10]), .B2(
        n2581), .ZN(n2760) );
  INV_X1 U2996 ( .A(n2586), .ZN(n485) );
  AOI222_X1 U2997 ( .A1(n2710), .A2(C21_DATA3_27), .B1(n2709), .B2(
        operand_ra_i[27]), .C1(dividend_q[27]), .C2(n2967), .ZN(n2586) );
  NAND2_X1 U2998 ( .A1(n2987), .A2(n2765), .ZN(n428) );
  AOI21_X1 U2999 ( .B1(C22_DATA3_11), .B2(n2571), .A(n2764), .ZN(n2765) );
  OAI21_X1 U3000 ( .B1(n2799), .B2(n92), .A(n2763), .ZN(n2764) );
  AOI22_X1 U3001 ( .A1(n2581), .A2(dividend_q[11]), .B1(result_o[11]), .B2(
        n2580), .ZN(n2763) );
  INV_X1 U3002 ( .A(n2585), .ZN(n484) );
  AOI222_X1 U3003 ( .A1(n2710), .A2(C21_DATA3_28), .B1(n2709), .B2(
        operand_ra_i[28]), .C1(dividend_q[28]), .C2(n2967), .ZN(n2585) );
  INV_X1 U3004 ( .A(n2711), .ZN(n483) );
  AOI222_X1 U3005 ( .A1(n2710), .A2(C21_DATA3_29), .B1(n2709), .B2(
        operand_ra_i[29]), .C1(dividend_q[29]), .C2(n2577), .ZN(n2711) );
  NAND2_X1 U3006 ( .A1(n2986), .A2(n2768), .ZN(n430) );
  AOI21_X1 U3007 ( .B1(C22_DATA3_13), .B2(n2571), .A(n2767), .ZN(n2768) );
  OAI21_X1 U3008 ( .B1(n2799), .B2(n90), .A(n2766), .ZN(n2767) );
  AOI22_X1 U3009 ( .A1(result_o[13]), .A2(n2580), .B1(dividend_q[13]), .B2(
        n2581), .ZN(n2766) );
  INV_X1 U3010 ( .A(n2584), .ZN(n482) );
  AOI222_X1 U3011 ( .A1(n2710), .A2(C21_DATA3_30), .B1(n2709), .B2(
        operand_ra_i[30]), .C1(dividend_q[30]), .C2(n2967), .ZN(n2584) );
  NAND2_X1 U3012 ( .A1(n2985), .A2(n2771), .ZN(n431) );
  AOI21_X1 U3013 ( .B1(C22_DATA3_14), .B2(n2571), .A(n2770), .ZN(n2771) );
  OAI21_X1 U3014 ( .B1(n2799), .B2(n8900), .A(n2769), .ZN(n2770) );
  AOI22_X1 U3015 ( .A1(n2581), .A2(dividend_q[14]), .B1(result_o[14]), .B2(
        n2580), .ZN(n2769) );
  NOR2_X1 U3016 ( .A1(n2573), .A2(n2524), .ZN(C1_Z_31) );
  NAND2_X1 U3017 ( .A1(n2574), .A2(divisor_q[31]), .ZN(n2615) );
  NOR2_X1 U3018 ( .A1(n2573), .A2(n2472), .ZN(C1_Z_0) );
  INV_X1 U3019 ( .A(operand_ra_i[0]), .ZN(n2707) );
  NOR2_X1 U3020 ( .A1(n2573), .A2(n2448), .ZN(C1_Z_1) );
  OAI21_X1 U3021 ( .B1(n2708), .B2(n2704), .A(n2705), .ZN(
        DP_OP_56J3_124_887_n102) );
  NAND2_X1 U3022 ( .A1(n2801), .A2(divisor_q[1]), .ZN(n2705) );
  NOR2_X1 U3023 ( .A1(n2573), .A2(n2447), .ZN(C1_Z_2) );
  OAI21_X1 U3024 ( .B1(n2567), .B2(n2701), .A(n2702), .ZN(
        DP_OP_56J3_124_887_n103) );
  NAND2_X1 U3025 ( .A1(n2801), .A2(divisor_q[2]), .ZN(n2702) );
  INV_X1 U3026 ( .A(operand_ra_i[2]), .ZN(n2701) );
  NOR2_X1 U3027 ( .A1(n2573), .A2(n2471), .ZN(C1_Z_3) );
  OAI21_X1 U3028 ( .B1(n2567), .B2(n2698), .A(n2699), .ZN(
        DP_OP_56J3_124_887_n104) );
  NAND2_X1 U3029 ( .A1(n2801), .A2(divisor_q[3]), .ZN(n2699) );
  INV_X1 U3030 ( .A(operand_ra_i[3]), .ZN(n2698) );
  NOR2_X1 U3031 ( .A1(n2573), .A2(n2481), .ZN(C1_Z_4) );
  OAI21_X1 U3032 ( .B1(n2567), .B2(n2695), .A(n2696), .ZN(
        DP_OP_56J3_124_887_n105) );
  NAND2_X1 U3033 ( .A1(n2801), .A2(divisor_q[4]), .ZN(n2696) );
  INV_X1 U3034 ( .A(operand_ra_i[4]), .ZN(n2695) );
  NOR2_X1 U3035 ( .A1(n2573), .A2(n2485), .ZN(C1_Z_5) );
  OAI21_X1 U3036 ( .B1(n2567), .B2(n2692), .A(n2693), .ZN(
        DP_OP_56J3_124_887_n106) );
  NAND2_X1 U3037 ( .A1(n2801), .A2(divisor_q[5]), .ZN(n2693) );
  INV_X1 U3038 ( .A(operand_ra_i[5]), .ZN(n2692) );
  NOR2_X1 U3039 ( .A1(n2573), .A2(n2482), .ZN(C1_Z_6) );
  OAI21_X1 U3040 ( .B1(n2567), .B2(n2689), .A(n2690), .ZN(
        DP_OP_56J3_124_887_n107) );
  NAND2_X1 U3041 ( .A1(n2801), .A2(divisor_q[6]), .ZN(n2690) );
  INV_X1 U3042 ( .A(operand_ra_i[6]), .ZN(n2689) );
  NOR2_X1 U3043 ( .A1(n2573), .A2(n2484), .ZN(C1_Z_7) );
  OAI21_X1 U3044 ( .B1(n2567), .B2(n2686), .A(n2687), .ZN(
        DP_OP_56J3_124_887_n108) );
  NAND2_X1 U3045 ( .A1(n2801), .A2(divisor_q[7]), .ZN(n2687) );
  INV_X1 U3046 ( .A(operand_ra_i[7]), .ZN(n2686) );
  NOR2_X1 U3047 ( .A1(n2573), .A2(n2478), .ZN(C1_Z_8) );
  OAI21_X1 U3048 ( .B1(n2566), .B2(n2683), .A(n2684), .ZN(
        DP_OP_56J3_124_887_n109) );
  NAND2_X1 U3049 ( .A1(n2801), .A2(divisor_q[8]), .ZN(n2684) );
  INV_X1 U3050 ( .A(operand_ra_i[8]), .ZN(n2683) );
  NOR2_X1 U3051 ( .A1(n2573), .A2(n2450), .ZN(C1_Z_9) );
  OAI21_X1 U3052 ( .B1(n2566), .B2(n2680), .A(n2681), .ZN(
        DP_OP_56J3_124_887_n110) );
  NAND2_X1 U3053 ( .A1(n2801), .A2(divisor_q[9]), .ZN(n2681) );
  INV_X1 U3054 ( .A(operand_ra_i[9]), .ZN(n2680) );
  NOR2_X1 U3055 ( .A1(n2573), .A2(n2476), .ZN(C1_Z_10) );
  OAI21_X1 U3056 ( .B1(n2566), .B2(n2677), .A(n2678), .ZN(
        DP_OP_56J3_124_887_n111) );
  NAND2_X1 U3057 ( .A1(n2574), .A2(divisor_q[10]), .ZN(n2678) );
  INV_X1 U3058 ( .A(operand_ra_i[10]), .ZN(n2677) );
  NOR2_X1 U3059 ( .A1(n2573), .A2(n2479), .ZN(C1_Z_11) );
  OAI21_X1 U3060 ( .B1(n2566), .B2(n2674), .A(n2675), .ZN(
        DP_OP_56J3_124_887_n112) );
  NAND2_X1 U3061 ( .A1(n2574), .A2(divisor_q[11]), .ZN(n2675) );
  INV_X1 U3062 ( .A(operand_ra_i[11]), .ZN(n2674) );
  NOR2_X1 U3063 ( .A1(n2573), .A2(n2477), .ZN(C1_Z_12) );
  OAI21_X1 U3064 ( .B1(n2566), .B2(n2671), .A(n2672), .ZN(
        DP_OP_56J3_124_887_n113) );
  NAND2_X1 U3065 ( .A1(n2574), .A2(divisor_q[12]), .ZN(n2672) );
  INV_X1 U3066 ( .A(operand_ra_i[12]), .ZN(n2671) );
  NOR2_X1 U3067 ( .A1(n2573), .A2(n2449), .ZN(C1_Z_13) );
  OAI21_X1 U3068 ( .B1(n2566), .B2(n2668), .A(n2669), .ZN(
        DP_OP_56J3_124_887_n114) );
  NAND2_X1 U3069 ( .A1(n2574), .A2(divisor_q[13]), .ZN(n2669) );
  INV_X1 U3070 ( .A(operand_ra_i[13]), .ZN(n2668) );
  NOR2_X1 U3071 ( .A1(n2573), .A2(n2480), .ZN(C1_Z_14) );
  OAI21_X1 U3072 ( .B1(n2566), .B2(n2665), .A(n2666), .ZN(
        DP_OP_56J3_124_887_n115) );
  NAND2_X1 U3073 ( .A1(n2574), .A2(divisor_q[14]), .ZN(n2666) );
  INV_X1 U3074 ( .A(operand_ra_i[14]), .ZN(n2665) );
  NOR2_X1 U3075 ( .A1(n2573), .A2(n2475), .ZN(C1_Z_15) );
  OAI21_X1 U3076 ( .B1(n2566), .B2(n2662), .A(n2663), .ZN(
        DP_OP_56J3_124_887_n116) );
  NAND2_X1 U3077 ( .A1(n2574), .A2(divisor_q[15]), .ZN(n2663) );
  INV_X1 U3078 ( .A(operand_ra_i[15]), .ZN(n2662) );
  NOR2_X1 U3079 ( .A1(n2573), .A2(n2493), .ZN(C1_Z_16) );
  OAI21_X1 U3080 ( .B1(n2566), .B2(n2659), .A(n2660), .ZN(
        DP_OP_56J3_124_887_n117) );
  NAND2_X1 U3081 ( .A1(n2574), .A2(divisor_q[16]), .ZN(n2660) );
  INV_X1 U3082 ( .A(operand_ra_i[16]), .ZN(n2659) );
  NOR2_X1 U3083 ( .A1(n2573), .A2(n2455), .ZN(C1_Z_17) );
  OAI21_X1 U3084 ( .B1(n2566), .B2(n2656), .A(n2657), .ZN(
        DP_OP_56J3_124_887_n118) );
  NAND2_X1 U3085 ( .A1(n2574), .A2(divisor_q[17]), .ZN(n2657) );
  INV_X1 U3086 ( .A(operand_ra_i[17]), .ZN(n2656) );
  NOR2_X1 U3087 ( .A1(n2573), .A2(n2491), .ZN(C1_Z_18) );
  OAI21_X1 U3088 ( .B1(n2566), .B2(n2653), .A(n2654), .ZN(
        DP_OP_56J3_124_887_n119) );
  NAND2_X1 U3089 ( .A1(n2574), .A2(divisor_q[18]), .ZN(n2654) );
  INV_X1 U3090 ( .A(operand_ra_i[18]), .ZN(n2653) );
  NOR2_X1 U3091 ( .A1(n2573), .A2(n2457), .ZN(C1_Z_19) );
  OAI21_X1 U3092 ( .B1(n2566), .B2(n2650), .A(n2651), .ZN(
        DP_OP_56J3_124_887_n120) );
  NAND2_X1 U3093 ( .A1(n2574), .A2(divisor_q[19]), .ZN(n2651) );
  INV_X1 U3094 ( .A(operand_ra_i[19]), .ZN(n2650) );
  NOR2_X1 U3095 ( .A1(n2573), .A2(n2497), .ZN(C1_Z_20) );
  OAI21_X1 U3096 ( .B1(n2566), .B2(n2647), .A(n2648), .ZN(
        DP_OP_56J3_124_887_n121) );
  NAND2_X1 U3097 ( .A1(n2574), .A2(divisor_q[20]), .ZN(n2648) );
  INV_X1 U3098 ( .A(operand_ra_i[20]), .ZN(n2647) );
  NOR2_X1 U3099 ( .A1(n2573), .A2(n2451), .ZN(C1_Z_21) );
  OAI21_X1 U3100 ( .B1(n2566), .B2(n2644), .A(n2645), .ZN(
        DP_OP_56J3_124_887_n122) );
  NAND2_X1 U3101 ( .A1(n2574), .A2(divisor_q[21]), .ZN(n2645) );
  INV_X1 U3102 ( .A(operand_ra_i[21]), .ZN(n2644) );
  NOR2_X1 U3103 ( .A1(n2573), .A2(n2490), .ZN(C1_Z_22) );
  OAI21_X1 U3104 ( .B1(n2566), .B2(n2641), .A(n2642), .ZN(
        DP_OP_56J3_124_887_n123) );
  NAND2_X1 U3105 ( .A1(n2574), .A2(divisor_q[22]), .ZN(n2642) );
  INV_X1 U3106 ( .A(operand_ra_i[22]), .ZN(n2641) );
  NOR2_X1 U3107 ( .A1(n2573), .A2(n2453), .ZN(C1_Z_23) );
  OAI21_X1 U3108 ( .B1(n2566), .B2(n2638), .A(n2639), .ZN(
        DP_OP_56J3_124_887_n124) );
  NAND2_X1 U3109 ( .A1(n2574), .A2(divisor_q[23]), .ZN(n2639) );
  INV_X1 U3110 ( .A(operand_ra_i[23]), .ZN(n2638) );
  NOR2_X1 U3111 ( .A1(n2573), .A2(n2498), .ZN(C1_Z_24) );
  OAI21_X1 U3112 ( .B1(n2566), .B2(n2635), .A(n2636), .ZN(
        DP_OP_56J3_124_887_n125) );
  NAND2_X1 U3113 ( .A1(n2574), .A2(divisor_q[24]), .ZN(n2636) );
  INV_X1 U3114 ( .A(operand_ra_i[24]), .ZN(n2635) );
  NOR2_X1 U3115 ( .A1(n2573), .A2(n2454), .ZN(C1_Z_25) );
  OAI21_X1 U3116 ( .B1(n2566), .B2(n2632), .A(n2633), .ZN(
        DP_OP_56J3_124_887_n126) );
  NAND2_X1 U3117 ( .A1(n2801), .A2(divisor_q[25]), .ZN(n2633) );
  INV_X1 U3118 ( .A(operand_ra_i[25]), .ZN(n2632) );
  NOR2_X1 U3119 ( .A1(n2573), .A2(n2489), .ZN(C1_Z_26) );
  OAI21_X1 U3120 ( .B1(n2566), .B2(n2629), .A(n2630), .ZN(
        DP_OP_56J3_124_887_n127) );
  NAND2_X1 U3121 ( .A1(n2801), .A2(divisor_q[26]), .ZN(n2630) );
  INV_X1 U3122 ( .A(operand_ra_i[26]), .ZN(n2629) );
  NOR2_X1 U3123 ( .A1(n2573), .A2(n2456), .ZN(C1_Z_27) );
  OAI21_X1 U3124 ( .B1(n2566), .B2(n2626), .A(n2627), .ZN(
        DP_OP_56J3_124_887_n128) );
  NAND2_X1 U3125 ( .A1(n2801), .A2(divisor_q[27]), .ZN(n2627) );
  INV_X1 U3126 ( .A(operand_ra_i[27]), .ZN(n2626) );
  NOR2_X1 U3127 ( .A1(n2573), .A2(n2496), .ZN(C1_Z_28) );
  OAI21_X1 U3128 ( .B1(n2566), .B2(n2623), .A(n2624), .ZN(
        DP_OP_56J3_124_887_n129) );
  NAND2_X1 U3129 ( .A1(n2801), .A2(divisor_q[28]), .ZN(n2624) );
  INV_X1 U3130 ( .A(operand_ra_i[28]), .ZN(n2623) );
  NOR2_X1 U3131 ( .A1(n2573), .A2(n2452), .ZN(C1_Z_29) );
  OAI21_X1 U3132 ( .B1(n2566), .B2(n2620), .A(n2621), .ZN(
        DP_OP_56J3_124_887_n130) );
  NAND2_X1 U3133 ( .A1(n2801), .A2(divisor_q[29]), .ZN(n2621) );
  INV_X1 U3134 ( .A(operand_ra_i[29]), .ZN(n2620) );
  NOR2_X1 U3135 ( .A1(n2573), .A2(n2492), .ZN(C1_Z_30) );
  OAI21_X1 U3136 ( .B1(n2566), .B2(n2617), .A(n2618), .ZN(
        DP_OP_56J3_124_887_n131) );
  NAND2_X1 U3137 ( .A1(n2574), .A2(divisor_q[30]), .ZN(n2618) );
  INV_X1 U3138 ( .A(operand_ra_i[30]), .ZN(n2617) );
  OAI21_X1 U3139 ( .B1(inst_rem_i), .B2(inst_div_i), .A(operand_ra_i[31]), 
        .ZN(n2583) );
  NOR3_X1 U3140 ( .A1(div_busy_q), .A2(rst_i), .A3(mul_busy_q), .ZN(n2582) );
  NAND2_X1 U3141 ( .A1(n2984), .A2(n2774), .ZN(n433) );
  AOI21_X1 U3142 ( .B1(C22_DATA3_16), .B2(n2571), .A(n2773), .ZN(n2774) );
  OAI21_X1 U3143 ( .B1(n2799), .B2(n87), .A(n2772), .ZN(n2773) );
  AOI22_X1 U3144 ( .A1(result_o[16]), .A2(n2580), .B1(dividend_q[16]), .B2(
        n2581), .ZN(n2772) );
  NAND2_X1 U3145 ( .A1(n2983), .A2(n2777), .ZN(n436) );
  AOI21_X1 U3146 ( .B1(C22_DATA3_19), .B2(n2571), .A(n2776), .ZN(n2777) );
  OAI21_X1 U3147 ( .B1(n2799), .B2(n8400), .A(n2775), .ZN(n2776) );
  AOI22_X1 U3148 ( .A1(n2581), .A2(dividend_q[19]), .B1(result_o[19]), .B2(
        n2580), .ZN(n2775) );
  NAND2_X1 U3149 ( .A1(n2982), .A2(n2780), .ZN(n437) );
  AOI21_X1 U3150 ( .B1(C22_DATA3_20), .B2(n2571), .A(n2779), .ZN(n2780) );
  OAI21_X1 U3151 ( .B1(n2799), .B2(n8300), .A(n2778), .ZN(n2779) );
  AOI22_X1 U3152 ( .A1(n2581), .A2(dividend_q[20]), .B1(result_o[20]), .B2(
        n2580), .ZN(n2778) );
  NAND2_X1 U3153 ( .A1(n2981), .A2(n2783), .ZN(n438) );
  AOI21_X1 U3154 ( .B1(C22_DATA3_21), .B2(n2571), .A(n2782), .ZN(n2783) );
  OAI21_X1 U3155 ( .B1(n2799), .B2(n8200), .A(n2781), .ZN(n2782) );
  AOI22_X1 U3156 ( .A1(result_o[21]), .A2(n2580), .B1(dividend_q[21]), .B2(
        n2581), .ZN(n2781) );
  NAND2_X1 U3157 ( .A1(n2980), .A2(n2786), .ZN(n439) );
  AOI21_X1 U3158 ( .B1(C22_DATA3_22), .B2(n2571), .A(n2785), .ZN(n2786) );
  OAI21_X1 U3159 ( .B1(n2799), .B2(n8100), .A(n2784), .ZN(n2785) );
  AOI22_X1 U3160 ( .A1(result_o[22]), .A2(n2580), .B1(dividend_q[22]), .B2(
        n2581), .ZN(n2784) );
  NAND2_X1 U3161 ( .A1(n2979), .A2(n2789), .ZN(n440) );
  AOI21_X1 U3162 ( .B1(C22_DATA3_23), .B2(n2571), .A(n2788), .ZN(n2789) );
  OAI21_X1 U3163 ( .B1(n2799), .B2(n8000), .A(n2787), .ZN(n2788) );
  AOI22_X1 U3164 ( .A1(result_o[23]), .A2(n2580), .B1(dividend_q[23]), .B2(
        n2581), .ZN(n2787) );
  NAND2_X1 U3165 ( .A1(n2978), .A2(n2792), .ZN(n441) );
  AOI21_X1 U3166 ( .B1(C22_DATA3_24), .B2(n2571), .A(n2791), .ZN(n2792) );
  OAI21_X1 U3167 ( .B1(n2799), .B2(n7900), .A(n2790), .ZN(n2791) );
  AOI22_X1 U3168 ( .A1(n2581), .A2(dividend_q[24]), .B1(result_o[24]), .B2(
        n2580), .ZN(n2790) );
  NAND2_X1 U3169 ( .A1(n2977), .A2(n2795), .ZN(n442) );
  AOI21_X1 U3170 ( .B1(C22_DATA3_25), .B2(n2571), .A(n2794), .ZN(n2795) );
  OAI21_X1 U3171 ( .B1(n2799), .B2(n7800), .A(n2793), .ZN(n2794) );
  AOI22_X1 U3172 ( .A1(result_o[25]), .A2(n2580), .B1(dividend_q[25]), .B2(
        n2581), .ZN(n2793) );
  AOI22_X1 U3173 ( .A1(n2581), .A2(dividend_q[28]), .B1(result_o[28]), .B2(
        n2580), .ZN(n2796) );
  OAI21_X1 U3174 ( .B1(n2799), .B2(n7400), .A(n2797), .ZN(n2798) );
  AOI22_X1 U3175 ( .A1(result_o[29]), .A2(n2580), .B1(dividend_q[29]), .B2(
        n2581), .ZN(n2797) );
  INV_X1 U3176 ( .A(n2976), .ZN(n2747) );
  AOI22_X1 U3177 ( .A1(n2570), .A2(quotient_q[0]), .B1(dividend_q[0]), .B2(
        n2569), .ZN(n2746) );
  NOR2_X1 U3178 ( .A1(div_inst_q), .A2(n104), .ZN(n2744) );
  AOI22_X1 U3179 ( .A1(n2570), .A2(quotient_q[7]), .B1(dividend_q[7]), .B2(
        n2569), .ZN(n2735) );
  AOI22_X1 U3180 ( .A1(n2570), .A2(quotient_q[6]), .B1(dividend_q[6]), .B2(
        n2569), .ZN(n2736) );
  AOI22_X1 U3181 ( .A1(n2570), .A2(quotient_q[5]), .B1(dividend_q[5]), .B2(
        n2569), .ZN(n2737) );
  AOI22_X1 U3182 ( .A1(n2570), .A2(quotient_q[4]), .B1(dividend_q[4]), .B2(
        n2569), .ZN(n2738) );
  AOI22_X1 U3183 ( .A1(n2570), .A2(quotient_q[3]), .B1(dividend_q[3]), .B2(
        n2569), .ZN(n2739) );
  AOI22_X1 U3184 ( .A1(n2570), .A2(quotient_q[2]), .B1(dividend_q[2]), .B2(
        n2569), .ZN(n2740) );
  AOI22_X1 U3185 ( .A1(n2570), .A2(quotient_q[1]), .B1(dividend_q[1]), .B2(
        n2569), .ZN(n2743) );
  AOI22_X1 U3186 ( .A1(n2745), .A2(quotient_q[11]), .B1(dividend_q[11]), .B2(
        n2569), .ZN(n2731) );
  AOI22_X1 U3187 ( .A1(n2570), .A2(quotient_q[10]), .B1(dividend_q[10]), .B2(
        n2569), .ZN(n2732) );
  AOI22_X1 U3188 ( .A1(n2570), .A2(quotient_q[9]), .B1(dividend_q[9]), .B2(
        n2569), .ZN(n2733) );
  AOI22_X1 U3189 ( .A1(n2570), .A2(quotient_q[8]), .B1(dividend_q[8]), .B2(
        n2569), .ZN(n2734) );
  NOR2_X1 U3190 ( .A1(n2483), .A2(n104), .ZN(n2745) );
  OR2_X1 U3191 ( .A1(mul_busy_q), .A2(n2973), .ZN(n2486) );
  OR2_X1 U3192 ( .A1(div_inst_q), .A2(n2976), .ZN(n2487) );
  AOI22_X1 U3193 ( .A1(n2570), .A2(quotient_q[30]), .B1(dividend_q[30]), .B2(
        n2569), .ZN(n2712) );
  AOI22_X1 U3194 ( .A1(n2745), .A2(quotient_q[29]), .B1(dividend_q[29]), .B2(
        n2569), .ZN(n2713) );
  AOI22_X1 U3195 ( .A1(n2745), .A2(quotient_q[26]), .B1(dividend_q[26]), .B2(
        n2569), .ZN(n2716) );
  AOI22_X1 U3196 ( .A1(n2745), .A2(quotient_q[25]), .B1(dividend_q[25]), .B2(
        n2569), .ZN(n2717) );
  AOI22_X1 U3197 ( .A1(n2745), .A2(quotient_q[28]), .B1(dividend_q[28]), .B2(
        n2569), .ZN(n2714) );
  AOI22_X1 U3198 ( .A1(n2745), .A2(quotient_q[27]), .B1(dividend_q[27]), .B2(
        n2569), .ZN(n2715) );
  AOI22_X1 U3199 ( .A1(n2745), .A2(quotient_q[24]), .B1(dividend_q[24]), .B2(
        n2569), .ZN(n2718) );
  AOI22_X1 U3200 ( .A1(n2745), .A2(quotient_q[23]), .B1(dividend_q[23]), .B2(
        n2744), .ZN(n2719) );
  AOI22_X1 U3201 ( .A1(n2745), .A2(quotient_q[22]), .B1(dividend_q[22]), .B2(
        n2744), .ZN(n2720) );
  AOI22_X1 U3202 ( .A1(n2745), .A2(quotient_q[21]), .B1(dividend_q[21]), .B2(
        n2744), .ZN(n2721) );
  AOI22_X1 U3203 ( .A1(n2745), .A2(quotient_q[20]), .B1(dividend_q[20]), .B2(
        n2744), .ZN(n2722) );
  AOI22_X1 U3204 ( .A1(n2570), .A2(quotient_q[19]), .B1(dividend_q[19]), .B2(
        n2744), .ZN(n2723) );
  AOI22_X1 U3205 ( .A1(n2570), .A2(quotient_q[18]), .B1(dividend_q[18]), .B2(
        n2744), .ZN(n2724) );
  AOI22_X1 U3206 ( .A1(n2570), .A2(quotient_q[17]), .B1(dividend_q[17]), .B2(
        n2744), .ZN(n2725) );
  AOI22_X1 U3207 ( .A1(n2570), .A2(quotient_q[16]), .B1(dividend_q[16]), .B2(
        n2744), .ZN(n2726) );
  AOI22_X1 U3208 ( .A1(n2570), .A2(quotient_q[15]), .B1(dividend_q[15]), .B2(
        n2744), .ZN(n2727) );
  AOI22_X1 U3209 ( .A1(n2570), .A2(quotient_q[14]), .B1(dividend_q[14]), .B2(
        n2744), .ZN(n2728) );
  AOI22_X1 U3210 ( .A1(n2570), .A2(quotient_q[13]), .B1(dividend_q[13]), .B2(
        n2744), .ZN(n2729) );
  AOI22_X1 U3211 ( .A1(n2570), .A2(quotient_q[12]), .B1(dividend_q[12]), .B2(
        n2744), .ZN(n2730) );
  AND2_X1 U3212 ( .A1(operand_ra_i[0]), .A2(n611), .ZN(n2529) );
  AND2_X1 U3213 ( .A1(operand_ra_i[1]), .A2(n611), .ZN(n2530) );
  AND2_X1 U3214 ( .A1(operand_ra_i[3]), .A2(n611), .ZN(n2531) );
  AND2_X1 U3215 ( .A1(operand_ra_i[4]), .A2(n611), .ZN(n2532) );
  AND2_X1 U3216 ( .A1(operand_ra_i[6]), .A2(n611), .ZN(n2533) );
  AND2_X1 U3217 ( .A1(operand_ra_i[7]), .A2(n611), .ZN(n2534) );
  INV_X1 U3218 ( .A(operand_rb_i[0]), .ZN(n2535) );
  AOI222_X1 U3219 ( .A1(n2710), .A2(C21_DATA3_2), .B1(n2709), .B2(
        operand_ra_i[2]), .C1(dividend_q[2]), .C2(n2577), .ZN(n2611) );
  INV_X1 U3220 ( .A(operand_rb_i[1]), .ZN(n2536) );
  AOI222_X1 U3221 ( .A1(n2710), .A2(C21_DATA3_1), .B1(n2709), .B2(
        operand_ra_i[1]), .C1(dividend_q[1]), .C2(n2577), .ZN(n2612) );
  INV_X1 U3222 ( .A(operand_ra_i[1]), .ZN(n2704) );
  XNOR2_X1 U3223 ( .A(sub_x_9_n1), .B(operand_rb_i[31]), .ZN(N200) );
  NOR4_X1 U3225 ( .A1(inst_mul_i), .A2(inst_mulhsu_i), .A3(inst_mulh_i), .A4(
        inst_mulhu_i), .ZN(n2804) );
  NAND2_X1 U3226 ( .A1(valid_i), .A2(n2802), .ZN(n2817) );
  NOR4_X1 U3227 ( .A1(q_mask_q[16]), .A2(q_mask_q[17]), .A3(q_mask_q[18]), 
        .A4(q_mask_q[19]), .ZN(n2814) );
  NOR4_X1 U3228 ( .A1(q_mask_q[15]), .A2(q_mask_q[20]), .A3(q_mask_q[21]), 
        .A4(q_mask_q[22]), .ZN(n2813) );
  NOR4_X1 U3229 ( .A1(q_mask_q[30]), .A2(q_mask_q[31]), .A3(q_mask_q[3]), .A4(
        q_mask_q[4]), .ZN(n2805) );
  NAND3_X1 U3230 ( .A1(n7100), .A2(n6400), .A3(n2805), .ZN(n2806) );
  NOR4_X1 U3231 ( .A1(q_mask_q[14]), .A2(q_mask_q[1]), .A3(n2473), .A4(n2806), 
        .ZN(n2812) );
  NOR4_X1 U3232 ( .A1(q_mask_q[23]), .A2(q_mask_q[24]), .A3(q_mask_q[25]), 
        .A4(q_mask_q[26]), .ZN(n2810) );
  NOR4_X1 U3233 ( .A1(q_mask_q[27]), .A2(q_mask_q[28]), .A3(q_mask_q[29]), 
        .A4(q_mask_q[2]), .ZN(n2809) );
  NOR4_X1 U3234 ( .A1(q_mask_q[5]), .A2(q_mask_q[6]), .A3(q_mask_q[8]), .A4(
        q_mask_q[9]), .ZN(n2808) );
  NOR4_X1 U3235 ( .A1(q_mask_q[10]), .A2(q_mask_q[11]), .A3(q_mask_q[12]), 
        .A4(q_mask_q[13]), .ZN(n2807) );
  AND4_X1 U3236 ( .A1(n2810), .A2(n2809), .A3(n2808), .A4(n2807), .ZN(n2811)
         );
  NAND4_X1 U3237 ( .A1(n2814), .A2(n2813), .A3(n2812), .A4(n2811), .ZN(n2972)
         );
  INV_X1 U3238 ( .A(n2817), .ZN(n2815) );
  OAI211_X1 U3239 ( .C1(inst_mulhsu_i), .C2(inst_mulh_i), .A(operand_ra_i[31]), 
        .B(n2815), .ZN(n402) );
  AND2_X1 U3240 ( .A1(operand_rb_i[0]), .A2(n611), .ZN(N56) );
  AND2_X1 U3241 ( .A1(operand_rb_i[1]), .A2(n611), .ZN(N57) );
  AOI21_X1 U3242 ( .B1(n2972), .B2(n2470), .A(rst_i), .ZN(N575) );
  AND2_X1 U3243 ( .A1(operand_rb_i[2]), .A2(n611), .ZN(N58) );
  AND2_X1 U3244 ( .A1(operand_rb_i[3]), .A2(n611), .ZN(N59) );
  AND2_X1 U3245 ( .A1(operand_rb_i[4]), .A2(n611), .ZN(N60) );
  AND2_X1 U3246 ( .A1(operand_rb_i[5]), .A2(n611), .ZN(N61) );
  AND2_X1 U3247 ( .A1(operand_rb_i[6]), .A2(n611), .ZN(N62) );
  AND2_X1 U3248 ( .A1(operand_rb_i[7]), .A2(n611), .ZN(N63) );
  AND2_X1 U3249 ( .A1(operand_rb_i[8]), .A2(n611), .ZN(N64) );
  AND2_X1 U3250 ( .A1(operand_rb_i[9]), .A2(n611), .ZN(N65) );
  AND2_X1 U3251 ( .A1(operand_rb_i[10]), .A2(n611), .ZN(N66) );
  AND2_X1 U3252 ( .A1(operand_rb_i[11]), .A2(n611), .ZN(N67) );
  AND2_X1 U3253 ( .A1(operand_rb_i[12]), .A2(n611), .ZN(N68) );
  AND2_X1 U3254 ( .A1(operand_rb_i[13]), .A2(n611), .ZN(N69) );
  AND2_X1 U3255 ( .A1(operand_rb_i[14]), .A2(n611), .ZN(N70) );
  AND2_X1 U3256 ( .A1(operand_rb_i[15]), .A2(n611), .ZN(N71) );
  AND2_X1 U3257 ( .A1(operand_rb_i[16]), .A2(n611), .ZN(N72) );
  AND2_X1 U3258 ( .A1(operand_rb_i[17]), .A2(n611), .ZN(N73) );
  AND2_X1 U3259 ( .A1(operand_rb_i[18]), .A2(n611), .ZN(N74) );
  AND2_X1 U3260 ( .A1(operand_rb_i[19]), .A2(n611), .ZN(N75) );
  AND2_X1 U3261 ( .A1(operand_rb_i[20]), .A2(n611), .ZN(N76) );
  AND2_X1 U3262 ( .A1(operand_rb_i[21]), .A2(n611), .ZN(N77) );
  AND2_X1 U3263 ( .A1(operand_rb_i[22]), .A2(n611), .ZN(N78) );
  AND2_X1 U3264 ( .A1(operand_rb_i[23]), .A2(n611), .ZN(N79) );
  AND2_X1 U3265 ( .A1(operand_rb_i[24]), .A2(n611), .ZN(N80) );
  AND2_X1 U3266 ( .A1(operand_rb_i[25]), .A2(n611), .ZN(N81) );
  AND2_X1 U3267 ( .A1(operand_rb_i[26]), .A2(n611), .ZN(N82) );
  AND2_X1 U3268 ( .A1(operand_rb_i[27]), .A2(n611), .ZN(N83) );
  AND2_X1 U3269 ( .A1(operand_rb_i[28]), .A2(n611), .ZN(N84) );
  AND2_X1 U3270 ( .A1(operand_rb_i[29]), .A2(n611), .ZN(N85) );
  AND2_X1 U3271 ( .A1(operand_rb_i[30]), .A2(n611), .ZN(N86) );
  INV_X1 U3272 ( .A(inst_mulh_i), .ZN(n2816) );
  NOR4_X1 U3273 ( .A1(inst_mulhsu_i), .A2(n2820), .A3(n2817), .A4(n2816), .ZN(
        N88) );
  NOR2_X1 U3274 ( .A1(inst_mul_i), .A2(n2499), .ZN(N89) );
  NOR2_X1 U3275 ( .A1(inst_divu_i), .A2(inst_remu_i), .ZN(n2818) );
  NOR2_X1 U3276 ( .A1(inst_div_i), .A2(inst_rem_i), .ZN(n2822) );
  OAI21_X1 U3277 ( .B1(n2511), .B2(n2572), .A(n2803), .ZN(n576) );
  NOR2_X1 U3278 ( .A1(n2822), .A2(n2820), .ZN(n2819) );
  NOR3_X1 U3279 ( .A1(n2822), .A2(n2821), .A3(n2820), .ZN(n2882) );
  AOI222_X1 U3280 ( .A1(divisor_q[62]), .A2(n406), .B1(operand_rb_i[31]), .B2(
        n2575), .C1(n2576), .C2(N200), .ZN(n386) );
  OAI22_X1 U3281 ( .A1(n7100), .A2(n2572), .B1(n2573), .B2(n2523), .ZN(n5750)
         );
  OAI22_X1 U3282 ( .A1(n2446), .A2(n2573), .B1(n2523), .B2(n2500), .ZN(n574)
         );
  OAI22_X1 U3283 ( .A1(n2446), .A2(n2572), .B1(n2464), .B2(n2573), .ZN(n573)
         );
  OAI22_X1 U3284 ( .A1(n2464), .A2(n2572), .B1(n2519), .B2(n2573), .ZN(n572)
         );
  OAI22_X1 U3285 ( .A1(n2458), .A2(n2573), .B1(n2519), .B2(n2500), .ZN(n571)
         );
  OAI22_X1 U3286 ( .A1(n2458), .A2(n2572), .B1(n2518), .B2(n2573), .ZN(n570)
         );
  OAI22_X1 U3287 ( .A1(n6400), .A2(n2573), .B1(n2518), .B2(n2500), .ZN(n569)
         );
  OAI22_X1 U3288 ( .A1(n6400), .A2(n2572), .B1(n2465), .B2(n2573), .ZN(n568)
         );
  OAI22_X1 U3289 ( .A1(n2465), .A2(n2572), .B1(n2520), .B2(n2573), .ZN(n567)
         );
  OAI22_X1 U3290 ( .A1(n2442), .A2(n2573), .B1(n2520), .B2(n2500), .ZN(n566)
         );
  OAI22_X1 U3291 ( .A1(n2442), .A2(n2572), .B1(n2462), .B2(n2573), .ZN(n565)
         );
  OAI22_X1 U3292 ( .A1(n2462), .A2(n2572), .B1(n2514), .B2(n2573), .ZN(n564)
         );
  OAI22_X1 U3293 ( .A1(n2514), .A2(n2572), .B1(n2469), .B2(n2573), .ZN(n563)
         );
  OAI22_X1 U3294 ( .A1(n2469), .A2(n2572), .B1(n2517), .B2(n2573), .ZN(n562)
         );
  OAI22_X1 U3295 ( .A1(n2443), .A2(n2573), .B1(n2517), .B2(n2572), .ZN(n561)
         );
  OAI22_X1 U3296 ( .A1(n2443), .A2(n2572), .B1(n2459), .B2(n2573), .ZN(n560)
         );
  OAI22_X1 U3297 ( .A1(n2459), .A2(n2572), .B1(n2512), .B2(n2573), .ZN(n559)
         );
  OAI22_X1 U3298 ( .A1(n2512), .A2(n2572), .B1(n2466), .B2(n2573), .ZN(n558)
         );
  OAI22_X1 U3299 ( .A1(n2466), .A2(n2572), .B1(n2521), .B2(n2573), .ZN(n557)
         );
  OAI22_X1 U3300 ( .A1(n2445), .A2(n2573), .B1(n2521), .B2(n2572), .ZN(n556)
         );
  OAI22_X1 U3301 ( .A1(n2445), .A2(n2572), .B1(n2467), .B2(n2573), .ZN(n555)
         );
  OAI22_X1 U3302 ( .A1(n2467), .A2(n2572), .B1(n2516), .B2(n2573), .ZN(n554)
         );
  OAI22_X1 U3303 ( .A1(n2516), .A2(n2572), .B1(n2460), .B2(n2573), .ZN(n553)
         );
  OAI22_X1 U3304 ( .A1(n2460), .A2(n2572), .B1(n2513), .B2(n2573), .ZN(n552)
         );
  OAI22_X1 U3305 ( .A1(n2513), .A2(n2572), .B1(n2468), .B2(n2573), .ZN(n551)
         );
  OAI22_X1 U3306 ( .A1(n2468), .A2(n2572), .B1(n2522), .B2(n2573), .ZN(n550)
         );
  OAI22_X1 U3307 ( .A1(n2444), .A2(n2573), .B1(n2522), .B2(n2500), .ZN(n549)
         );
  OAI22_X1 U3308 ( .A1(n2444), .A2(n2572), .B1(n2463), .B2(n2573), .ZN(n548)
         );
  OAI22_X1 U3309 ( .A1(n2463), .A2(n2572), .B1(n2515), .B2(n2573), .ZN(n547)
         );
  OAI22_X1 U3310 ( .A1(n2515), .A2(n2572), .B1(n2461), .B2(n2573), .ZN(n546)
         );
  OAI22_X1 U3311 ( .A1(n2461), .A2(n2572), .B1(n2511), .B2(n2573), .ZN(n545)
         );
  AOI22_X1 U3312 ( .A1(n2574), .A2(divisor_q[33]), .B1(operand_rb_i[1]), .B2(
        n2881), .ZN(n2824) );
  AOI22_X1 U3313 ( .A1(divisor_q[32]), .A2(n406), .B1(n2576), .B2(N170), .ZN(
        n2823) );
  NAND2_X1 U3314 ( .A1(n2824), .A2(n2823), .ZN(n543) );
  AOI22_X1 U3315 ( .A1(n2574), .A2(divisor_q[34]), .B1(operand_rb_i[2]), .B2(
        n2881), .ZN(n2826) );
  AOI22_X1 U3316 ( .A1(divisor_q[33]), .A2(n406), .B1(n2882), .B2(N171), .ZN(
        n2825) );
  NAND2_X1 U3317 ( .A1(n2826), .A2(n2825), .ZN(n542) );
  AOI22_X1 U3318 ( .A1(n2574), .A2(divisor_q[35]), .B1(operand_rb_i[3]), .B2(
        n2881), .ZN(n2828) );
  AOI22_X1 U3319 ( .A1(divisor_q[34]), .A2(n406), .B1(n2576), .B2(N172), .ZN(
        n2827) );
  NAND2_X1 U3320 ( .A1(n2828), .A2(n2827), .ZN(n541) );
  AOI22_X1 U3321 ( .A1(n2574), .A2(divisor_q[36]), .B1(operand_rb_i[4]), .B2(
        n2575), .ZN(n2830) );
  AOI22_X1 U3322 ( .A1(divisor_q[35]), .A2(n406), .B1(n2576), .B2(N173), .ZN(
        n2829) );
  NAND2_X1 U3323 ( .A1(n2830), .A2(n2829), .ZN(n540) );
  AOI22_X1 U3324 ( .A1(n2574), .A2(divisor_q[37]), .B1(operand_rb_i[5]), .B2(
        n2575), .ZN(n2832) );
  AOI22_X1 U3325 ( .A1(divisor_q[36]), .A2(n406), .B1(n2576), .B2(N174), .ZN(
        n2831) );
  NAND2_X1 U3326 ( .A1(n2832), .A2(n2831), .ZN(n539) );
  AOI22_X1 U3327 ( .A1(n2574), .A2(divisor_q[38]), .B1(operand_rb_i[6]), .B2(
        n2881), .ZN(n2834) );
  AOI22_X1 U3328 ( .A1(divisor_q[37]), .A2(n406), .B1(n2576), .B2(N175), .ZN(
        n2833) );
  NAND2_X1 U3329 ( .A1(n2834), .A2(n2833), .ZN(n538) );
  AOI22_X1 U3330 ( .A1(n2574), .A2(divisor_q[39]), .B1(operand_rb_i[7]), .B2(
        n2881), .ZN(n2836) );
  AOI22_X1 U3331 ( .A1(divisor_q[38]), .A2(n406), .B1(n2576), .B2(N176), .ZN(
        n2835) );
  NAND2_X1 U3332 ( .A1(n2836), .A2(n2835), .ZN(n537) );
  AOI22_X1 U3333 ( .A1(n2574), .A2(divisor_q[40]), .B1(operand_rb_i[8]), .B2(
        n2881), .ZN(n2838) );
  AOI22_X1 U3334 ( .A1(divisor_q[39]), .A2(n406), .B1(n2576), .B2(N177), .ZN(
        n2837) );
  NAND2_X1 U3335 ( .A1(n2838), .A2(n2837), .ZN(n536) );
  AOI22_X1 U3336 ( .A1(n2801), .A2(divisor_q[41]), .B1(operand_rb_i[9]), .B2(
        n2881), .ZN(n2840) );
  AOI22_X1 U3337 ( .A1(divisor_q[40]), .A2(n406), .B1(n2576), .B2(N178), .ZN(
        n2839) );
  NAND2_X1 U3338 ( .A1(n2840), .A2(n2839), .ZN(n535) );
  AOI22_X1 U3339 ( .A1(n2574), .A2(divisor_q[42]), .B1(operand_rb_i[10]), .B2(
        n2881), .ZN(n2842) );
  AOI22_X1 U3340 ( .A1(divisor_q[41]), .A2(n406), .B1(n2576), .B2(N179), .ZN(
        n2841) );
  NAND2_X1 U3341 ( .A1(n2842), .A2(n2841), .ZN(n534) );
  AOI22_X1 U3342 ( .A1(n2801), .A2(divisor_q[43]), .B1(operand_rb_i[11]), .B2(
        n2881), .ZN(n2844) );
  AOI22_X1 U3343 ( .A1(divisor_q[42]), .A2(n406), .B1(n2576), .B2(N180), .ZN(
        n2843) );
  NAND2_X1 U3344 ( .A1(n2844), .A2(n2843), .ZN(n533) );
  AOI22_X1 U3345 ( .A1(n2801), .A2(divisor_q[44]), .B1(operand_rb_i[12]), .B2(
        n2881), .ZN(n2846) );
  AOI22_X1 U3346 ( .A1(divisor_q[43]), .A2(n406), .B1(n2576), .B2(N181), .ZN(
        n2845) );
  NAND2_X1 U3347 ( .A1(n2846), .A2(n2845), .ZN(n532) );
  AOI22_X1 U3348 ( .A1(n2574), .A2(divisor_q[45]), .B1(operand_rb_i[13]), .B2(
        n2881), .ZN(n2848) );
  AOI22_X1 U3349 ( .A1(divisor_q[44]), .A2(n406), .B1(n2576), .B2(N182), .ZN(
        n2847) );
  NAND2_X1 U3350 ( .A1(n2848), .A2(n2847), .ZN(n531) );
  AOI22_X1 U3351 ( .A1(n2801), .A2(divisor_q[46]), .B1(operand_rb_i[14]), .B2(
        n2575), .ZN(n2850) );
  AOI22_X1 U3352 ( .A1(divisor_q[45]), .A2(n406), .B1(n2576), .B2(N183), .ZN(
        n2849) );
  NAND2_X1 U3353 ( .A1(n2850), .A2(n2849), .ZN(n530) );
  AOI22_X1 U3354 ( .A1(n2801), .A2(divisor_q[47]), .B1(operand_rb_i[15]), .B2(
        n2575), .ZN(n2852) );
  AOI22_X1 U3355 ( .A1(divisor_q[46]), .A2(n406), .B1(n2576), .B2(N184), .ZN(
        n2851) );
  NAND2_X1 U3356 ( .A1(n2852), .A2(n2851), .ZN(n529) );
  AOI22_X1 U3357 ( .A1(n2801), .A2(divisor_q[48]), .B1(operand_rb_i[16]), .B2(
        n2575), .ZN(n2854) );
  AOI22_X1 U3358 ( .A1(divisor_q[47]), .A2(n406), .B1(n2576), .B2(N185), .ZN(
        n2853) );
  NAND2_X1 U3359 ( .A1(n2854), .A2(n2853), .ZN(n528) );
  AOI22_X1 U3360 ( .A1(n2574), .A2(divisor_q[49]), .B1(operand_rb_i[17]), .B2(
        n2575), .ZN(n2856) );
  AOI22_X1 U3361 ( .A1(divisor_q[48]), .A2(n406), .B1(n2576), .B2(N186), .ZN(
        n2855) );
  NAND2_X1 U3362 ( .A1(n2856), .A2(n2855), .ZN(n527) );
  AOI22_X1 U3363 ( .A1(n2801), .A2(divisor_q[50]), .B1(operand_rb_i[18]), .B2(
        n2881), .ZN(n2858) );
  AOI22_X1 U3364 ( .A1(divisor_q[49]), .A2(n406), .B1(n2576), .B2(N187), .ZN(
        n2857) );
  NAND2_X1 U3365 ( .A1(n2858), .A2(n2857), .ZN(n526) );
  AOI22_X1 U3366 ( .A1(n2574), .A2(divisor_q[51]), .B1(operand_rb_i[19]), .B2(
        n2575), .ZN(n2860) );
  AOI22_X1 U3367 ( .A1(divisor_q[50]), .A2(n406), .B1(n2882), .B2(N188), .ZN(
        n2859) );
  NAND2_X1 U3368 ( .A1(n2860), .A2(n2859), .ZN(n525) );
  AOI22_X1 U3369 ( .A1(n2574), .A2(divisor_q[52]), .B1(operand_rb_i[20]), .B2(
        n2575), .ZN(n2862) );
  AOI22_X1 U3370 ( .A1(divisor_q[51]), .A2(n406), .B1(n2882), .B2(N189), .ZN(
        n2861) );
  NAND2_X1 U3371 ( .A1(n2862), .A2(n2861), .ZN(n524) );
  AOI22_X1 U3372 ( .A1(n2801), .A2(divisor_q[53]), .B1(operand_rb_i[21]), .B2(
        n2575), .ZN(n2864) );
  AOI22_X1 U3373 ( .A1(divisor_q[52]), .A2(n406), .B1(n2882), .B2(N190), .ZN(
        n2863) );
  NAND2_X1 U3374 ( .A1(n2864), .A2(n2863), .ZN(n523) );
  AOI22_X1 U3375 ( .A1(n2574), .A2(divisor_q[54]), .B1(operand_rb_i[22]), .B2(
        n2575), .ZN(n2866) );
  AOI22_X1 U3376 ( .A1(divisor_q[53]), .A2(n406), .B1(n2576), .B2(N191), .ZN(
        n2865) );
  NAND2_X1 U3377 ( .A1(n2866), .A2(n2865), .ZN(n522) );
  AOI22_X1 U3378 ( .A1(n2574), .A2(divisor_q[55]), .B1(operand_rb_i[23]), .B2(
        n2575), .ZN(n2868) );
  AOI22_X1 U3379 ( .A1(divisor_q[54]), .A2(n406), .B1(n2576), .B2(N192), .ZN(
        n2867) );
  NAND2_X1 U3380 ( .A1(n2868), .A2(n2867), .ZN(n521) );
  AOI22_X1 U3381 ( .A1(n2574), .A2(divisor_q[56]), .B1(operand_rb_i[24]), .B2(
        n2575), .ZN(n2870) );
  AOI22_X1 U3382 ( .A1(divisor_q[55]), .A2(n406), .B1(n2882), .B2(N193), .ZN(
        n2869) );
  NAND2_X1 U3383 ( .A1(n2870), .A2(n2869), .ZN(n520) );
  AOI22_X1 U3384 ( .A1(n2574), .A2(divisor_q[57]), .B1(operand_rb_i[25]), .B2(
        n2575), .ZN(n2872) );
  AOI22_X1 U3385 ( .A1(divisor_q[56]), .A2(n406), .B1(n2576), .B2(N194), .ZN(
        n2871) );
  NAND2_X1 U3386 ( .A1(n2872), .A2(n2871), .ZN(n519) );
  AOI22_X1 U3387 ( .A1(n2574), .A2(divisor_q[58]), .B1(operand_rb_i[26]), .B2(
        n2575), .ZN(n2874) );
  AOI22_X1 U3388 ( .A1(divisor_q[57]), .A2(n406), .B1(n2576), .B2(N195), .ZN(
        n2873) );
  NAND2_X1 U3389 ( .A1(n2874), .A2(n2873), .ZN(n518) );
  AOI22_X1 U3390 ( .A1(n2574), .A2(divisor_q[59]), .B1(operand_rb_i[27]), .B2(
        n2575), .ZN(n2876) );
  AOI22_X1 U3391 ( .A1(divisor_q[58]), .A2(n406), .B1(n2576), .B2(N196), .ZN(
        n2875) );
  NAND2_X1 U3392 ( .A1(n2876), .A2(n2875), .ZN(n517) );
  AOI22_X1 U3393 ( .A1(n2574), .A2(divisor_q[60]), .B1(operand_rb_i[28]), .B2(
        n2575), .ZN(n2878) );
  AOI22_X1 U3394 ( .A1(divisor_q[59]), .A2(n406), .B1(n2882), .B2(N197), .ZN(
        n2877) );
  NAND2_X1 U3395 ( .A1(n2878), .A2(n2877), .ZN(n516) );
  AOI22_X1 U3396 ( .A1(n2574), .A2(divisor_q[61]), .B1(operand_rb_i[29]), .B2(
        n2575), .ZN(n2880) );
  AOI22_X1 U3397 ( .A1(divisor_q[60]), .A2(n406), .B1(n2882), .B2(N198), .ZN(
        n2879) );
  NAND2_X1 U3398 ( .A1(n2880), .A2(n2879), .ZN(n515) );
  AOI22_X1 U3399 ( .A1(n2574), .A2(divisor_q[62]), .B1(operand_rb_i[30]), .B2(
        n2575), .ZN(n2884) );
  AOI22_X1 U3400 ( .A1(divisor_q[61]), .A2(n406), .B1(n2576), .B2(N199), .ZN(
        n2883) );
  NAND2_X1 U3401 ( .A1(n2884), .A2(n2883), .ZN(n514) );
  OAI21_X1 U3402 ( .B1(n2452), .B2(divisor_q[29]), .A(n2496), .ZN(n2885) );
  INV_X1 U3403 ( .A(n2885), .ZN(n2886) );
  AOI22_X1 U3404 ( .A1(n2886), .A2(divisor_q[28]), .B1(divisor_q[29]), .B2(
        n2452), .ZN(n2889) );
  OAI22_X1 U3405 ( .A1(divisor_q[31]), .A2(n2524), .B1(divisor_q[30]), .B2(
        n2492), .ZN(n2954) );
  NOR4_X1 U3406 ( .A1(divisor_q[34]), .A2(divisor_q[35]), .A3(divisor_q[46]), 
        .A4(divisor_q[36]), .ZN(n2888) );
  NOR4_X1 U3407 ( .A1(divisor_q[37]), .A2(divisor_q[47]), .A3(divisor_q[48]), 
        .A4(divisor_q[49]), .ZN(n2887) );
  OAI211_X1 U3408 ( .C1(n2889), .C2(n2954), .A(n2888), .B(n2887), .ZN(n2965)
         );
  NOR4_X1 U3409 ( .A1(divisor_q[55]), .A2(divisor_q[53]), .A3(divisor_q[54]), 
        .A4(divisor_q[56]), .ZN(n2963) );
  AOI21_X1 U3410 ( .B1(divisor_q[31]), .B2(n2524), .A(divisor_q[52]), .ZN(
        n2962) );
  OAI211_X1 U3411 ( .C1(n2524), .C2(divisor_q[31]), .A(n2492), .B(
        divisor_q[30]), .ZN(n2890) );
  INV_X1 U3412 ( .A(n2890), .ZN(n2896) );
  NOR4_X1 U3413 ( .A1(divisor_q[62]), .A2(divisor_q[60]), .A3(divisor_q[32]), 
        .A4(divisor_q[33]), .ZN(n2894) );
  NOR4_X1 U3414 ( .A1(divisor_q[57]), .A2(divisor_q[58]), .A3(divisor_q[59]), 
        .A4(divisor_q[61]), .ZN(n2893) );
  NOR4_X1 U3415 ( .A1(divisor_q[42]), .A2(divisor_q[43]), .A3(divisor_q[44]), 
        .A4(divisor_q[45]), .ZN(n2892) );
  NOR4_X1 U3416 ( .A1(divisor_q[38]), .A2(divisor_q[41]), .A3(divisor_q[39]), 
        .A4(divisor_q[40]), .ZN(n2891) );
  NAND4_X1 U3417 ( .A1(n2894), .A2(n2893), .A3(n2892), .A4(n2891), .ZN(n2895)
         );
  NOR4_X1 U3418 ( .A1(n2896), .A2(divisor_q[50]), .A3(divisor_q[51]), .A4(
        n2895), .ZN(n2961) );
  OAI211_X1 U3419 ( .C1(divisor_q[27]), .C2(n2456), .A(divisor_q[26]), .B(
        n2489), .ZN(n2901) );
  OAI211_X1 U3420 ( .C1(n2454), .C2(divisor_q[25]), .A(n2498), .B(
        divisor_q[24]), .ZN(n2897) );
  INV_X1 U3421 ( .A(n2897), .ZN(n2899) );
  OAI22_X1 U3422 ( .A1(n2456), .A2(divisor_q[27]), .B1(n2489), .B2(
        divisor_q[26]), .ZN(n2902) );
  INV_X1 U3423 ( .A(n2902), .ZN(n2898) );
  OAI221_X1 U3424 ( .B1(n2899), .B2(divisor_q[25]), .C1(n2899), .C2(n2454), 
        .A(n2898), .ZN(n2900) );
  OAI211_X1 U3425 ( .C1(dividend_q[27]), .C2(n2502), .A(n2901), .B(n2900), 
        .ZN(n2959) );
  NOR2_X1 U3426 ( .A1(divisor_q[25]), .A2(n2454), .ZN(n2903) );
  AOI211_X1 U3427 ( .C1(dividend_q[24]), .C2(n2507), .A(n2903), .B(n2902), 
        .ZN(n2958) );
  OAI21_X1 U3428 ( .B1(n2451), .B2(divisor_q[21]), .A(n2497), .ZN(n2904) );
  INV_X1 U3429 ( .A(n2904), .ZN(n2905) );
  AOI22_X1 U3430 ( .A1(n2905), .A2(divisor_q[20]), .B1(divisor_q[21]), .B2(
        n2451), .ZN(n2953) );
  OAI22_X1 U3431 ( .A1(divisor_q[23]), .A2(n2453), .B1(divisor_q[22]), .B2(
        n2490), .ZN(n2952) );
  OAI21_X1 U3432 ( .B1(n2453), .B2(divisor_q[23]), .A(n2490), .ZN(n2906) );
  INV_X1 U3433 ( .A(n2906), .ZN(n2907) );
  AOI22_X1 U3434 ( .A1(n2907), .A2(divisor_q[22]), .B1(divisor_q[23]), .B2(
        n2453), .ZN(n2951) );
  NOR2_X1 U3435 ( .A1(divisor_q[11]), .A2(n2479), .ZN(n2913) );
  OAI22_X1 U3436 ( .A1(n2450), .A2(divisor_q[9]), .B1(n2476), .B2(
        divisor_q[10]), .ZN(n2912) );
  INV_X1 U3437 ( .A(n2912), .ZN(n2910) );
  AOI22_X1 U3438 ( .A1(n2478), .A2(divisor_q[8]), .B1(n2450), .B2(divisor_q[9]), .ZN(n2908) );
  INV_X1 U3439 ( .A(n2908), .ZN(n2909) );
  AOI22_X1 U3440 ( .A1(n2910), .A2(n2909), .B1(divisor_q[10]), .B2(n2476), 
        .ZN(n2911) );
  OAI22_X1 U3441 ( .A1(n2913), .A2(n2911), .B1(dividend_q[11]), .B2(n2508), 
        .ZN(n2930) );
  AOI211_X1 U3442 ( .C1(dividend_q[8]), .C2(n2504), .A(n2913), .B(n2912), .ZN(
        n2929) );
  AOI22_X1 U3443 ( .A1(divisor_q[3]), .A2(n2471), .B1(divisor_q[2]), .B2(n2447), .ZN(n2917) );
  OAI21_X1 U3444 ( .B1(divisor_q[1]), .B2(n2448), .A(divisor_q[0]), .ZN(n2914)
         );
  OAI22_X1 U3445 ( .A1(dividend_q[0]), .A2(n2914), .B1(dividend_q[1]), .B2(
        n2510), .ZN(n2915) );
  OAI21_X1 U3446 ( .B1(divisor_q[2]), .B2(n2447), .A(n2915), .ZN(n2916) );
  AOI22_X1 U3447 ( .A1(dividend_q[3]), .A2(n2503), .B1(n2917), .B2(n2916), 
        .ZN(n2920) );
  AND2_X1 U3448 ( .A1(divisor_q[4]), .A2(n2481), .ZN(n2919) );
  NAND2_X1 U3449 ( .A1(dividend_q[5]), .A2(n2494), .ZN(n2918) );
  OAI221_X1 U3450 ( .B1(divisor_q[4]), .B2(n2481), .C1(n2920), .C2(n2919), .A(
        n2918), .ZN(n2921) );
  OAI21_X1 U3451 ( .B1(dividend_q[5]), .B2(n2494), .A(n2921), .ZN(n2924) );
  AND2_X1 U3452 ( .A1(divisor_q[6]), .A2(n2482), .ZN(n2923) );
  NAND2_X1 U3453 ( .A1(dividend_q[7]), .A2(n2495), .ZN(n2922) );
  OAI221_X1 U3454 ( .B1(divisor_q[6]), .B2(n2482), .C1(n2924), .C2(n2923), .A(
        n2922), .ZN(n2925) );
  OAI21_X1 U3455 ( .B1(dividend_q[7]), .B2(n2495), .A(n2925), .ZN(n2928) );
  NOR2_X1 U3456 ( .A1(divisor_q[14]), .A2(n2480), .ZN(n2934) );
  OAI22_X1 U3457 ( .A1(divisor_q[13]), .A2(n2449), .B1(divisor_q[12]), .B2(
        n2477), .ZN(n2926) );
  AOI211_X1 U3458 ( .C1(dividend_q[15]), .C2(n2488), .A(n2934), .B(n2926), 
        .ZN(n2927) );
  OAI221_X1 U3459 ( .B1(n2930), .B2(n2929), .C1(n2930), .C2(n2928), .A(n2927), 
        .ZN(n2939) );
  NAND2_X1 U3460 ( .A1(dividend_q[15]), .A2(n2488), .ZN(n2936) );
  OAI21_X1 U3461 ( .B1(n2449), .B2(divisor_q[13]), .A(n2477), .ZN(n2931) );
  INV_X1 U3462 ( .A(n2931), .ZN(n2932) );
  AOI22_X1 U3463 ( .A1(n2932), .A2(divisor_q[12]), .B1(divisor_q[13]), .B2(
        n2449), .ZN(n2933) );
  OAI22_X1 U3464 ( .A1(n2934), .A2(n2933), .B1(dividend_q[14]), .B2(n2509), 
        .ZN(n2935) );
  AOI22_X1 U3465 ( .A1(divisor_q[15]), .A2(n2475), .B1(n2936), .B2(n2935), 
        .ZN(n2938) );
  OAI22_X1 U3466 ( .A1(divisor_q[19]), .A2(n2457), .B1(divisor_q[18]), .B2(
        n2491), .ZN(n2941) );
  OAI22_X1 U3467 ( .A1(divisor_q[17]), .A2(n2455), .B1(divisor_q[16]), .B2(
        n2493), .ZN(n2937) );
  AOI211_X1 U3468 ( .C1(n2939), .C2(n2938), .A(n2941), .B(n2937), .ZN(n2949)
         );
  OAI211_X1 U3469 ( .C1(divisor_q[19]), .C2(n2457), .A(divisor_q[18]), .B(
        n2491), .ZN(n2945) );
  OAI211_X1 U3470 ( .C1(n2455), .C2(divisor_q[17]), .A(n2493), .B(
        divisor_q[16]), .ZN(n2940) );
  INV_X1 U3471 ( .A(n2940), .ZN(n2943) );
  INV_X1 U3472 ( .A(n2941), .ZN(n2942) );
  OAI221_X1 U3473 ( .B1(n2943), .B2(divisor_q[17]), .C1(n2943), .C2(n2455), 
        .A(n2942), .ZN(n2944) );
  OAI211_X1 U3474 ( .C1(dividend_q[19]), .C2(n2501), .A(n2945), .B(n2944), 
        .ZN(n2948) );
  NOR2_X1 U3475 ( .A1(divisor_q[21]), .A2(n2451), .ZN(n2946) );
  AOI211_X1 U3476 ( .C1(dividend_q[20]), .C2(n2505), .A(n2946), .B(n2952), 
        .ZN(n2947) );
  OAI21_X1 U3477 ( .B1(n2949), .B2(n2948), .A(n2947), .ZN(n2950) );
  OAI211_X1 U3478 ( .C1(n2953), .C2(n2952), .A(n2951), .B(n2950), .ZN(n2957)
         );
  NOR2_X1 U3479 ( .A1(divisor_q[29]), .A2(n2452), .ZN(n2955) );
  AOI211_X1 U3480 ( .C1(dividend_q[28]), .C2(n2506), .A(n2955), .B(n2954), 
        .ZN(n2956) );
  OAI221_X1 U3481 ( .B1(n2959), .B2(n2958), .C1(n2959), .C2(n2957), .A(n2956), 
        .ZN(n2960) );
  NAND4_X1 U3482 ( .A1(n2963), .A2(n2962), .A3(n2961), .A4(n2960), .ZN(n2964)
         );
  OAI21_X1 U3483 ( .B1(n2965), .B2(n2964), .A(n2968), .ZN(n2966) );
  NAND2_X1 U3484 ( .A1(n2966), .A2(n2500), .ZN(n2967) );
  OAI21_X1 U3485 ( .B1(inst_divu_i), .B2(inst_div_i), .A(n2969), .ZN(n2970) );
  NOR2_X1 U3486 ( .A1(rst_i), .A2(n2972), .ZN(n2974) );
  NAND2_X1 U3487 ( .A1(n2974), .A2(n104), .ZN(n2976) );
  INV_X1 U3488 ( .A(n2974), .ZN(n2975) );
  AOI22_X1 U3489 ( .A1(n2579), .A2(mult_result_w[25]), .B1(mult_result_w[57]), 
        .B2(n2993), .ZN(n2977) );
  AOI22_X1 U3490 ( .A1(n2579), .A2(mult_result_w[24]), .B1(n2993), .B2(
        mult_result_w[56]), .ZN(n2978) );
  AOI22_X1 U3491 ( .A1(n2579), .A2(mult_result_w[23]), .B1(n2993), .B2(
        mult_result_w[55]), .ZN(n2979) );
  AOI22_X1 U3492 ( .A1(n2579), .A2(mult_result_w[22]), .B1(n2993), .B2(
        mult_result_w[54]), .ZN(n2980) );
  AOI22_X1 U3493 ( .A1(n2579), .A2(mult_result_w[21]), .B1(n2993), .B2(
        mult_result_w[53]), .ZN(n2981) );
  AOI22_X1 U3494 ( .A1(n2579), .A2(mult_result_w[20]), .B1(n2993), .B2(
        mult_result_w[52]), .ZN(n2982) );
  AOI22_X1 U3495 ( .A1(n2579), .A2(mult_result_w[19]), .B1(n2578), .B2(
        mult_result_w[51]), .ZN(n2983) );
  AOI22_X1 U3496 ( .A1(n2579), .A2(mult_result_w[16]), .B1(n2578), .B2(
        mult_result_w[48]), .ZN(n2984) );
  AOI22_X1 U3497 ( .A1(n2579), .A2(mult_result_w[14]), .B1(n2578), .B2(
        mult_result_w[46]), .ZN(n2985) );
  AOI22_X1 U3498 ( .A1(n2579), .A2(mult_result_w[13]), .B1(n2578), .B2(
        mult_result_w[45]), .ZN(n2986) );
  AOI22_X1 U3499 ( .A1(n2579), .A2(mult_result_w[11]), .B1(n2578), .B2(
        mult_result_w[43]), .ZN(n2987) );
  AOI22_X1 U3500 ( .A1(n2579), .A2(mult_result_w[10]), .B1(n2578), .B2(
        mult_result_w[42]), .ZN(n2988) );
  AOI22_X1 U3501 ( .A1(n2579), .A2(mult_result_w[7]), .B1(n2578), .B2(
        mult_result_w[39]), .ZN(n2989) );
  AOI22_X1 U3502 ( .A1(n2994), .A2(mult_result_w[6]), .B1(n2578), .B2(
        mult_result_w[38]), .ZN(n2990) );
  AOI22_X1 U3503 ( .A1(n2994), .A2(mult_result_w[4]), .B1(n2578), .B2(
        mult_result_w[36]), .ZN(n2991) );
  AOI22_X1 U3504 ( .A1(n2994), .A2(mult_result_w[3]), .B1(n2578), .B2(
        mult_result_w[35]), .ZN(n2992) );
endmodule


module riscv_core ( clk_i, rst_i, intr_i, reset_vector_i, cpu_id_i, mem_i_rd_o, 
        mem_i_pc_o, mem_i_accept_i, mem_i_valid_i, mem_i_inst_i, mem_i_flush_o, 
        mem_i_invalidate_o, mem_i_error_i, mem_d_addr_o, mem_d_data_wr_o, 
        mem_d_rd_o, mem_d_wr_o, mem_d_data_rd_i, mem_d_accept_i, mem_d_ack_i, 
        mem_d_cacheable_o, mem_d_req_tag_o, mem_d_invalidate_o, 
        mem_d_writeback_o, mem_d_flush_o, mem_d_error_i, mem_d_resp_tag_i );
  input [31:0] reset_vector_i;
  input [31:0] cpu_id_i;
  output [31:0] mem_i_pc_o;
  input [31:0] mem_i_inst_i;
  output [31:0] mem_d_addr_o;
  output [31:0] mem_d_data_wr_o;
  output [3:0] mem_d_wr_o;
  input [31:0] mem_d_data_rd_i;
  output [10:0] mem_d_req_tag_o;
  input [10:0] mem_d_resp_tag_i;
  input clk_i, rst_i, intr_i, mem_i_accept_i, mem_i_valid_i, mem_i_error_i,
         mem_d_accept_i, mem_d_ack_i, mem_d_error_i;
  output mem_i_rd_o, mem_i_flush_o, mem_i_invalidate_o, mem_d_rd_o,
         mem_d_cacheable_o, mem_d_invalidate_o, mem_d_writeback_o,
         mem_d_flush_o;
  wire   rd_wr_en_q, state_q_0_, muldiv_ready_w, exception_w, inst_mul_w,
         inst_mulh_w, inst_mulhsu_w, inst_mulhu_w, inst_div_w, inst_divu_w,
         inst_rem_w, inst_remu_w, invalid_inst_r, mem_misaligned_w,
         n_0_net__29_, n_0_net__27_, n_0_net__25_, n_0_net__23_, n_0_net__17_,
         n_0_net__13_, n_0_net__4_, n_1_net_, u_branch_N127, u_branch_N125,
         u_branch_N120, u_lsu_N16, u_lsu_N14, n57, n143, n144, n145, n146,
         n147, n154, n155, n156, n157, n158, n159, n160, n161, n162, n1370,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1463, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2872,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2919, C1_Z_2, U4_RSOP_173_C3_DATA1_30,
         U4_RSOP_173_C3_DATA1_29, U4_RSOP_173_C3_DATA1_28,
         U4_RSOP_173_C3_DATA1_27, U4_RSOP_173_C3_DATA1_26,
         U4_RSOP_173_C3_DATA1_25, U4_RSOP_173_C3_DATA1_24,
         U4_RSOP_173_C3_DATA1_23, U4_RSOP_173_C3_DATA1_22,
         U4_RSOP_173_C3_DATA1_21, U4_RSOP_173_C3_DATA1_20,
         U4_RSOP_173_C3_DATA1_19, U4_RSOP_173_C3_DATA1_17,
         U4_RSOP_173_C3_DATA1_16, U4_RSOP_173_C3_DATA1_15,
         U4_RSOP_173_C3_DATA1_13, U4_RSOP_173_C3_DATA1_12,
         U4_RSOP_173_C3_DATA1_11, U4_RSOP_173_C3_DATA1_8,
         U4_RSOP_173_C3_DATA1_7, U4_RSOP_173_C3_DATA1_4,
         U4_RSOP_173_C3_DATA1_3, U4_RSOP_173_C3_DATA1_0, add_x_67_B_4_,
         add_x_67_B_3_, add_x_67_B_1_, add_x_67_n32, add_x_67_n31,
         add_x_67_n30, add_x_67_n29, add_x_67_n28, add_x_67_n27, add_x_67_n26,
         add_x_67_n25, add_x_67_n24, add_x_67_n23, add_x_67_n22, add_x_67_n21,
         add_x_67_n20, add_x_67_n19, add_x_67_n18, add_x_67_n17, add_x_67_n16,
         add_x_67_n15, add_x_67_n14, add_x_67_n13, add_x_67_n12, add_x_67_n11,
         add_x_67_n10, add_x_67_n9, add_x_67_n8, add_x_67_n7, add_x_67_n6,
         add_x_67_n5, add_x_67_n4, add_x_67_n3, add_x_67_n2, sub_x_59_n94,
         sub_x_59_n93, sub_x_59_n92, sub_x_59_n85, sub_x_59_n84, sub_x_59_n78,
         sub_x_59_n77, sub_x_59_n76, sub_x_59_n65, sub_x_59_n63, sub_x_59_n59,
         sub_x_59_n41, sub_x_59_n39, sub_x_59_n29, sub_x_59_n28, sub_x_59_n17,
         sub_x_59_n8, sub_x_59_n7, sub_x_59_n1, sub_x_60_n94, sub_x_60_n93,
         sub_x_60_n92, sub_x_60_n84, sub_x_60_n78, sub_x_60_n77, sub_x_60_n76,
         sub_x_60_n61, sub_x_60_n29, sub_x_60_n28, sub_x_60_n12, sub_x_60_n11,
         sub_x_60_n9, sub_x_60_n8, sub_x_60_n1, DP_OP_181_135_5161_n121,
         DP_OP_181_135_5161_n120, DP_OP_181_135_5161_n119,
         DP_OP_181_135_5161_n118, DP_OP_181_135_5161_n117,
         DP_OP_181_135_5161_n116, DP_OP_181_135_5161_n115,
         DP_OP_181_135_5161_n114, DP_OP_181_135_5161_n113,
         DP_OP_181_135_5161_n112, DP_OP_181_135_5161_n111,
         DP_OP_181_135_5161_n110, DP_OP_181_135_5161_n109,
         DP_OP_181_135_5161_n108, DP_OP_181_135_5161_n107,
         DP_OP_181_135_5161_n106, DP_OP_181_135_5161_n105,
         DP_OP_181_135_5161_n104, DP_OP_181_135_5161_n103,
         DP_OP_181_135_5161_n102, DP_OP_181_135_5161_n100,
         DP_OP_181_135_5161_n99, DP_OP_181_135_5161_n98,
         DP_OP_181_135_5161_n97, DP_OP_181_135_5161_n96,
         DP_OP_181_135_5161_n95, DP_OP_181_135_5161_n94,
         DP_OP_181_135_5161_n93, DP_OP_181_135_5161_n92,
         DP_OP_181_135_5161_n91, DP_OP_181_135_5161_n89,
         DP_OP_181_135_5161_n88, DP_OP_181_135_5161_n87,
         DP_OP_181_135_5161_n86, DP_OP_181_135_5161_n85,
         DP_OP_181_135_5161_n84, DP_OP_181_135_5161_n83,
         DP_OP_181_135_5161_n82, DP_OP_181_135_5161_n81,
         DP_OP_181_135_5161_n79, DP_OP_181_135_5161_n78,
         DP_OP_181_135_5161_n77, DP_OP_181_135_5161_n76,
         DP_OP_181_135_5161_n75, DP_OP_181_135_5161_n74,
         DP_OP_181_135_5161_n73, DP_OP_181_135_5161_n72,
         DP_OP_181_135_5161_n70, DP_OP_181_135_5161_n32,
         DP_OP_181_135_5161_n30, DP_OP_181_135_5161_n29,
         DP_OP_181_135_5161_n28, DP_OP_181_135_5161_n26,
         DP_OP_181_135_5161_n25, DP_OP_181_135_5161_n24,
         DP_OP_181_135_5161_n22, DP_OP_181_135_5161_n21,
         DP_OP_181_135_5161_n20, DP_OP_181_135_5161_n18,
         DP_OP_181_135_5161_n17, DP_OP_181_135_5161_n16,
         DP_OP_181_135_5161_n14, DP_OP_181_135_5161_n13,
         DP_OP_181_135_5161_n12, DP_OP_181_135_5161_n11,
         DP_OP_181_135_5161_n10, DP_OP_181_135_5161_n9, DP_OP_181_135_5161_n8,
         DP_OP_181_135_5161_n7, DP_OP_181_135_5161_n5, DP_OP_181_135_5161_n4,
         DP_OP_181_135_5161_n3, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38;
  wire   [31:0] alu_a_q;
  wire   [31:0] alu_b_q;
  wire   [1023:0] reg_file;
  wire   [31:0] rs1_val_gpr_w;
  wire   [31:0] rs2_val_gpr_w;
  wire   [31:0] csr_data_w;
  wire   [31:0] muldiv_result_w;
  wire   [31:0] csr_mepc_w;
  wire   [31:0] mem_addr_w;
  assign mem_i_flush_o = 1'b0;
  assign mem_i_invalidate_o = 1'b0;
  assign mem_d_cacheable_o = 1'b0;
  assign mem_d_req_tag_o[10] = 1'b0;
  assign mem_d_req_tag_o[9] = 1'b0;
  assign mem_d_req_tag_o[8] = 1'b0;
  assign mem_d_req_tag_o[7] = 1'b0;
  assign mem_d_req_tag_o[6] = 1'b0;
  assign mem_d_req_tag_o[5] = 1'b0;
  assign mem_d_req_tag_o[4] = 1'b0;
  assign mem_d_req_tag_o[3] = 1'b0;
  assign mem_d_req_tag_o[2] = 1'b0;
  assign mem_d_req_tag_o[1] = 1'b0;
  assign mem_d_req_tag_o[0] = 1'b0;
  assign mem_d_invalidate_o = 1'b0;
  assign mem_d_writeback_o = 1'b0;
  assign mem_d_flush_o = 1'b0;
  assign mem_d_addr_o[0] = 1'b0;
  assign mem_d_addr_o[1] = 1'b0;

  uriscv_csr_SUPPORT_CSR1_SUPPORT_MCYCLE1_SUPPORT_MTIMECMP0_SUPPORT_MSCRATCH0_SUPPORT_MIP_MIE0_SUPPORT_MTVEC0_SUPPORT_MTVAL0_SUPPORT_MULDIV1 u_csr ( 
        .clk_i(clk_i), .rst_i(rst_i), .intr_i(intr_i), .isr_vector_i({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cpu_id_i(cpu_id_i), 
        .valid_i(mem_i_valid_i), .pc_i(mem_i_pc_o), .opcode_i({
        mem_i_inst_i[31:2], 1'b0, 1'b0}), .rs1_val_i({rs1_val_gpr_w[31:8], 
        n3523, rs1_val_gpr_w[6:4], n3524, rs1_val_gpr_w[2:1], n3521}), 
        .rs2_val_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .csr_rdata_o(csr_data_w), .excpn_invalid_inst_i(invalid_inst_r), 
        .excpn_lsu_align_i(mem_misaligned_w), .mem_addr_i({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .csr_mepc_o(csr_mepc_w), .exception_o(
        exception_w), .exception_type_o({SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6}), .exception_pc_o({
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38}) );
  uriscv_muldiv genblk1_u_muldiv ( .clk_i(clk_i), .rst_i(rst_i), .valid_i(
        n_1_net_), .inst_mul_i(inst_mul_w), .inst_mulh_i(inst_mulh_w), 
        .inst_mulhsu_i(inst_mulhsu_w), .inst_mulhu_i(inst_mulhu_w), 
        .inst_div_i(inst_div_w), .inst_divu_i(inst_divu_w), .inst_rem_i(
        inst_rem_w), .inst_remu_i(inst_remu_w), .operand_ra_i({
        rs1_val_gpr_w[31:8], n3523, rs1_val_gpr_w[6:4], n3524, 
        rs1_val_gpr_w[2:1], n3521}), .operand_rb_i(rs2_val_gpr_w), .ready_o(
        muldiv_ready_w), .result_o(muldiv_result_w) );
  DFF_X1 pc_q_reg_0_ ( .D(n2916), .CK(clk_i), .Q(mem_i_pc_o[0]), .QN(n3801) );
  DFF_X1 state_q_reg_1_ ( .D(n2917), .CK(clk_i), .Q(n3837), .QN(n57) );
  DFF_X1 state_q_reg_0_ ( .D(n2919), .CK(clk_i), .Q(state_q_0_) );
  DFF_X1 rd_wr_en_q_reg ( .D(n2875), .CK(clk_i), .Q(rd_wr_en_q) );
  DFF_X1 rd_q_reg_4_ ( .D(n2880), .CK(clk_i), .QN(n143) );
  DFF_X1 pc_q_reg_1_ ( .D(n2915), .CK(clk_i), .Q(mem_i_pc_o[1]) );
  DFF_X1 pc_q_reg_2_ ( .D(n2914), .CK(clk_i), .Q(mem_i_pc_o[2]), .QN(n3771) );
  DFF_X1 pc_q_reg_3_ ( .D(n2913), .CK(clk_i), .Q(mem_i_pc_o[3]), .QN(n3823) );
  DFF_X1 pc_q_reg_4_ ( .D(n2912), .CK(clk_i), .Q(mem_i_pc_o[4]), .QN(n3824) );
  DFF_X1 pc_q_reg_5_ ( .D(n2911), .CK(clk_i), .Q(mem_i_pc_o[5]), .QN(n3828) );
  DFF_X1 pc_q_reg_6_ ( .D(n2910), .CK(clk_i), .Q(mem_i_pc_o[6]), .QN(n3827) );
  DFF_X1 pc_q_reg_7_ ( .D(n2909), .CK(clk_i), .Q(mem_i_pc_o[7]), .QN(n3826) );
  DFF_X1 pc_q_reg_8_ ( .D(n2908), .CK(clk_i), .Q(mem_i_pc_o[8]), .QN(n3825) );
  DFF_X1 pc_q_reg_9_ ( .D(n2907), .CK(clk_i), .Q(mem_i_pc_o[9]), .QN(n3822) );
  DFF_X1 pc_q_reg_10_ ( .D(n2906), .CK(clk_i), .Q(mem_i_pc_o[10]), .QN(n3821)
         );
  DFF_X1 pc_q_reg_11_ ( .D(n2905), .CK(clk_i), .Q(mem_i_pc_o[11]), .QN(n3820)
         );
  DFF_X1 pc_q_reg_12_ ( .D(n2904), .CK(clk_i), .Q(mem_i_pc_o[12]), .QN(n3819)
         );
  DFF_X1 pc_q_reg_13_ ( .D(n2903), .CK(clk_i), .Q(mem_i_pc_o[13]), .QN(n3818)
         );
  DFF_X1 pc_q_reg_14_ ( .D(n2902), .CK(clk_i), .Q(mem_i_pc_o[14]), .QN(n3817)
         );
  DFF_X1 pc_q_reg_15_ ( .D(n2901), .CK(clk_i), .Q(mem_i_pc_o[15]), .QN(n3816)
         );
  DFF_X1 pc_q_reg_16_ ( .D(n2900), .CK(clk_i), .Q(mem_i_pc_o[16]), .QN(n3863)
         );
  DFF_X1 pc_q_reg_17_ ( .D(n2899), .CK(clk_i), .Q(mem_i_pc_o[17]), .QN(n3862)
         );
  DFF_X1 pc_q_reg_18_ ( .D(n2898), .CK(clk_i), .Q(mem_i_pc_o[18]), .QN(n3861)
         );
  DFF_X1 pc_q_reg_19_ ( .D(n2897), .CK(clk_i), .Q(mem_i_pc_o[19]), .QN(n3860)
         );
  DFF_X1 pc_q_reg_20_ ( .D(n2896), .CK(clk_i), .Q(mem_i_pc_o[20]), .QN(n3859)
         );
  DFF_X1 pc_q_reg_21_ ( .D(n2895), .CK(clk_i), .Q(mem_i_pc_o[21]), .QN(n3858)
         );
  DFF_X1 pc_q_reg_22_ ( .D(n2894), .CK(clk_i), .Q(mem_i_pc_o[22]), .QN(n3857)
         );
  DFF_X1 pc_q_reg_23_ ( .D(n2893), .CK(clk_i), .Q(mem_i_pc_o[23]), .QN(n3856)
         );
  DFF_X1 pc_q_reg_24_ ( .D(n2892), .CK(clk_i), .Q(mem_i_pc_o[24]), .QN(n3855)
         );
  DFF_X1 pc_q_reg_25_ ( .D(n2891), .CK(clk_i), .Q(mem_i_pc_o[25]), .QN(n3854)
         );
  DFF_X1 pc_q_reg_26_ ( .D(n2890), .CK(clk_i), .Q(mem_i_pc_o[26]), .QN(n3853)
         );
  DFF_X1 pc_q_reg_27_ ( .D(n2889), .CK(clk_i), .Q(mem_i_pc_o[27]), .QN(n3852)
         );
  DFF_X1 pc_q_reg_28_ ( .D(n2888), .CK(clk_i), .Q(mem_i_pc_o[28]), .QN(n3872)
         );
  DFF_X1 pc_q_reg_31_ ( .D(n2885), .CK(clk_i), .Q(mem_i_pc_o[31]), .QN(n3869)
         );
  DFF_X1 alu_b_q_reg_25_ ( .D(n2849), .CK(clk_i), .Q(alu_b_q[25]) );
  DFF_X1 alu_b_q_reg_30_ ( .D(n2844), .CK(clk_i), .Q(alu_b_q[30]) );
  DFF_X1 mem_rd_q_reg ( .D(n1463), .CK(clk_i), .QN(mem_d_rd_o) );
  DFF_X1 mem_addr_q_reg_31_ ( .D(n1461), .CK(clk_i), .QN(mem_d_addr_o[31]) );
  DFF_X1 mem_addr_q_reg_30_ ( .D(n1460), .CK(clk_i), .QN(mem_d_addr_o[30]) );
  DFF_X1 mem_addr_q_reg_29_ ( .D(n1459), .CK(clk_i), .QN(mem_d_addr_o[29]) );
  DFF_X1 mem_addr_q_reg_28_ ( .D(n1458), .CK(clk_i), .QN(mem_d_addr_o[28]) );
  DFF_X1 mem_addr_q_reg_27_ ( .D(n1457), .CK(clk_i), .QN(mem_d_addr_o[27]) );
  DFF_X1 mem_addr_q_reg_26_ ( .D(n1456), .CK(clk_i), .QN(mem_d_addr_o[26]) );
  DFF_X1 mem_addr_q_reg_25_ ( .D(n1455), .CK(clk_i), .QN(mem_d_addr_o[25]) );
  DFF_X1 mem_addr_q_reg_24_ ( .D(n1454), .CK(clk_i), .QN(mem_d_addr_o[24]) );
  DFF_X1 mem_addr_q_reg_23_ ( .D(n1453), .CK(clk_i), .QN(mem_d_addr_o[23]) );
  DFF_X1 mem_addr_q_reg_22_ ( .D(n1452), .CK(clk_i), .QN(mem_d_addr_o[22]) );
  DFF_X1 mem_addr_q_reg_21_ ( .D(n1451), .CK(clk_i), .QN(mem_d_addr_o[21]) );
  DFF_X1 mem_addr_q_reg_20_ ( .D(n1450), .CK(clk_i), .QN(mem_d_addr_o[20]) );
  DFF_X1 mem_addr_q_reg_19_ ( .D(n1449), .CK(clk_i), .QN(mem_d_addr_o[19]) );
  DFF_X1 mem_addr_q_reg_18_ ( .D(n1448), .CK(clk_i), .QN(mem_d_addr_o[18]) );
  DFF_X1 mem_addr_q_reg_17_ ( .D(n1447), .CK(clk_i), .QN(mem_d_addr_o[17]) );
  DFF_X1 mem_addr_q_reg_16_ ( .D(n1446), .CK(clk_i), .QN(mem_d_addr_o[16]) );
  DFF_X1 mem_addr_q_reg_15_ ( .D(n1445), .CK(clk_i), .QN(mem_d_addr_o[15]) );
  DFF_X1 mem_addr_q_reg_14_ ( .D(n1444), .CK(clk_i), .QN(mem_d_addr_o[14]) );
  DFF_X1 mem_addr_q_reg_13_ ( .D(n1443), .CK(clk_i), .QN(mem_d_addr_o[13]) );
  DFF_X1 mem_addr_q_reg_12_ ( .D(n1442), .CK(clk_i), .QN(mem_d_addr_o[12]) );
  DFF_X1 mem_addr_q_reg_11_ ( .D(n1441), .CK(clk_i), .QN(mem_d_addr_o[11]) );
  DFF_X1 mem_addr_q_reg_10_ ( .D(n1440), .CK(clk_i), .QN(mem_d_addr_o[10]) );
  DFF_X1 mem_addr_q_reg_9_ ( .D(n1439), .CK(clk_i), .QN(mem_d_addr_o[9]) );
  DFF_X1 mem_addr_q_reg_8_ ( .D(n1438), .CK(clk_i), .QN(mem_d_addr_o[8]) );
  DFF_X1 mem_addr_q_reg_7_ ( .D(n1437), .CK(clk_i), .QN(mem_d_addr_o[7]) );
  DFF_X1 mem_addr_q_reg_6_ ( .D(n1436), .CK(clk_i), .QN(mem_d_addr_o[6]) );
  DFF_X1 mem_addr_q_reg_5_ ( .D(n1435), .CK(clk_i), .QN(mem_d_addr_o[5]) );
  DFF_X1 mem_addr_q_reg_4_ ( .D(n1434), .CK(clk_i), .QN(mem_d_addr_o[4]) );
  DFF_X1 mem_addr_q_reg_3_ ( .D(n1433), .CK(clk_i), .QN(mem_d_addr_o[3]) );
  DFF_X1 mem_addr_q_reg_2_ ( .D(n1432), .CK(clk_i), .QN(mem_d_addr_o[2]) );
  DFF_X1 mem_data_q_reg_31_ ( .D(n2842), .CK(clk_i), .Q(mem_d_data_wr_o[31])
         );
  DFF_X1 mem_data_q_reg_30_ ( .D(n2841), .CK(clk_i), .Q(mem_d_data_wr_o[30])
         );
  DFF_X1 mem_data_q_reg_29_ ( .D(n2840), .CK(clk_i), .Q(mem_d_data_wr_o[29])
         );
  DFF_X1 mem_data_q_reg_28_ ( .D(n2839), .CK(clk_i), .Q(mem_d_data_wr_o[28])
         );
  DFF_X1 mem_data_q_reg_27_ ( .D(n2838), .CK(clk_i), .Q(mem_d_data_wr_o[27])
         );
  DFF_X1 mem_data_q_reg_26_ ( .D(n2837), .CK(clk_i), .Q(mem_d_data_wr_o[26])
         );
  DFF_X1 mem_data_q_reg_25_ ( .D(n2836), .CK(clk_i), .Q(mem_d_data_wr_o[25])
         );
  DFF_X1 mem_data_q_reg_24_ ( .D(n2835), .CK(clk_i), .Q(mem_d_data_wr_o[24])
         );
  DFF_X1 mem_data_q_reg_23_ ( .D(n2834), .CK(clk_i), .Q(mem_d_data_wr_o[23])
         );
  DFF_X1 mem_data_q_reg_22_ ( .D(n2833), .CK(clk_i), .Q(mem_d_data_wr_o[22])
         );
  DFF_X1 mem_data_q_reg_21_ ( .D(n2832), .CK(clk_i), .Q(mem_d_data_wr_o[21])
         );
  DFF_X1 mem_data_q_reg_20_ ( .D(n2831), .CK(clk_i), .Q(mem_d_data_wr_o[20])
         );
  DFF_X1 mem_data_q_reg_19_ ( .D(n2830), .CK(clk_i), .Q(mem_d_data_wr_o[19])
         );
  DFF_X1 mem_data_q_reg_18_ ( .D(n2829), .CK(clk_i), .Q(mem_d_data_wr_o[18])
         );
  DFF_X1 mem_data_q_reg_17_ ( .D(n2828), .CK(clk_i), .Q(mem_d_data_wr_o[17])
         );
  DFF_X1 mem_data_q_reg_16_ ( .D(n2827), .CK(clk_i), .Q(mem_d_data_wr_o[16])
         );
  DFF_X1 mem_data_q_reg_15_ ( .D(n2826), .CK(clk_i), .Q(mem_d_data_wr_o[15])
         );
  DFF_X1 mem_data_q_reg_14_ ( .D(n2825), .CK(clk_i), .Q(mem_d_data_wr_o[14])
         );
  DFF_X1 mem_data_q_reg_13_ ( .D(n2824), .CK(clk_i), .Q(mem_d_data_wr_o[13])
         );
  DFF_X1 mem_data_q_reg_12_ ( .D(n2823), .CK(clk_i), .Q(mem_d_data_wr_o[12])
         );
  DFF_X1 mem_data_q_reg_11_ ( .D(n2822), .CK(clk_i), .Q(mem_d_data_wr_o[11])
         );
  DFF_X1 mem_data_q_reg_10_ ( .D(n2821), .CK(clk_i), .Q(mem_d_data_wr_o[10])
         );
  DFF_X1 mem_data_q_reg_9_ ( .D(n2820), .CK(clk_i), .Q(mem_d_data_wr_o[9]) );
  DFF_X1 mem_data_q_reg_8_ ( .D(n2819), .CK(clk_i), .Q(mem_d_data_wr_o[8]) );
  DFF_X1 mem_data_q_reg_7_ ( .D(n1387), .CK(clk_i), .QN(mem_d_data_wr_o[7]) );
  DFF_X1 mem_data_q_reg_6_ ( .D(n1386), .CK(clk_i), .QN(mem_d_data_wr_o[6]) );
  DFF_X1 mem_data_q_reg_5_ ( .D(n1385), .CK(clk_i), .QN(mem_d_data_wr_o[5]) );
  DFF_X1 mem_data_q_reg_4_ ( .D(n1384), .CK(clk_i), .QN(mem_d_data_wr_o[4]) );
  DFF_X1 mem_data_q_reg_3_ ( .D(n1383), .CK(clk_i), .QN(mem_d_data_wr_o[3]) );
  DFF_X1 mem_data_q_reg_2_ ( .D(n1382), .CK(clk_i), .QN(mem_d_data_wr_o[2]) );
  DFF_X1 mem_data_q_reg_1_ ( .D(n1381), .CK(clk_i), .QN(mem_d_data_wr_o[1]) );
  DFF_X1 mem_data_q_reg_0_ ( .D(n1380), .CK(clk_i), .QN(mem_d_data_wr_o[0]) );
  DFF_X1 mem_wr_q_reg_3_ ( .D(n2818), .CK(clk_i), .Q(mem_d_wr_o[3]) );
  DFF_X1 mem_wr_q_reg_2_ ( .D(n2817), .CK(clk_i), .Q(mem_d_wr_o[2]) );
  DFF_X1 mem_wr_q_reg_1_ ( .D(n2816), .CK(clk_i), .Q(mem_d_wr_o[1]), .QN(n4708) );
  DFF_X1 mem_wr_q_reg_0_ ( .D(n1370), .CK(clk_i), .QN(mem_d_wr_o[0]) );
  DFF_X1 load_half_q_reg ( .D(n2814), .CK(clk_i), .QN(n159) );
  DFF_X1 alu_a_q_reg_7_ ( .D(n2803), .CK(clk_i), .Q(alu_a_q[7]) );
  DFF_X1 alu_a_q_reg_14_ ( .D(n2796), .CK(clk_i), .Q(alu_a_q[14]) );
  DFF_X1 alu_a_q_reg_10_ ( .D(n2800), .CK(clk_i), .Q(alu_a_q[10]) );
  DFF_X1 reg_file_reg_31__31_ ( .D(n1787), .CK(clk_i), .Q(reg_file[31]), .QN(
        n4707) );
  DFF_X1 reg_file_reg_30__31_ ( .D(n1788), .CK(clk_i), .Q(reg_file[63]), .QN(
        n4183) );
  DFF_X1 reg_file_reg_29__31_ ( .D(n1789), .CK(clk_i), .Q(reg_file[95]), .QN(
        n4182) );
  DFF_X1 reg_file_reg_28__31_ ( .D(n1790), .CK(clk_i), .Q(reg_file[127]), .QN(
        n4706) );
  DFF_X1 reg_file_reg_27__31_ ( .D(n1791), .CK(clk_i), .Q(reg_file[159]), .QN(
        n4395) );
  DFF_X1 reg_file_reg_26__31_ ( .D(n1792), .CK(clk_i), .Q(reg_file[191]), .QN(
        n4394) );
  DFF_X1 reg_file_reg_25__31_ ( .D(n1793), .CK(clk_i), .Q(reg_file[223]), .QN(
        n4393) );
  DFF_X1 reg_file_reg_24__31_ ( .D(n1794), .CK(clk_i), .Q(reg_file[255]), .QN(
        n4699) );
  DFF_X1 reg_file_reg_23__31_ ( .D(n1795), .CK(clk_i), .Q(reg_file[287]), .QN(
        n4705) );
  DFF_X1 reg_file_reg_22__31_ ( .D(n1796), .CK(clk_i), .Q(reg_file[319]), .QN(
        n4181) );
  DFF_X1 reg_file_reg_21__31_ ( .D(n1797), .CK(clk_i), .Q(reg_file[351]), .QN(
        n4180) );
  DFF_X1 reg_file_reg_20__31_ ( .D(n1798), .CK(clk_i), .Q(reg_file[383]), .QN(
        n4704) );
  DFF_X1 reg_file_reg_19__31_ ( .D(n1799), .CK(clk_i), .Q(reg_file[415]), .QN(
        n4392) );
  DFF_X1 reg_file_reg_18__31_ ( .D(n1800), .CK(clk_i), .Q(reg_file[447]), .QN(
        n4391) );
  DFF_X1 reg_file_reg_17__31_ ( .D(n1801), .CK(clk_i), .Q(reg_file[479]), .QN(
        n4390) );
  DFF_X1 reg_file_reg_16__31_ ( .D(n1802), .CK(clk_i), .Q(reg_file[511]), .QN(
        n4698) );
  DFF_X1 reg_file_reg_15__31_ ( .D(n1803), .CK(clk_i), .Q(reg_file[543]), .QN(
        n4703) );
  DFF_X1 reg_file_reg_14__31_ ( .D(n1804), .CK(clk_i), .Q(reg_file[575]), .QN(
        n4179) );
  DFF_X1 reg_file_reg_13__31_ ( .D(n1805), .CK(clk_i), .Q(reg_file[607]), .QN(
        n4178) );
  DFF_X1 reg_file_reg_12__31_ ( .D(n1806), .CK(clk_i), .Q(reg_file[639]), .QN(
        n4702) );
  DFF_X1 reg_file_reg_11__31_ ( .D(n1807), .CK(clk_i), .Q(reg_file[671]), .QN(
        n4389) );
  DFF_X1 reg_file_reg_10__31_ ( .D(n1808), .CK(clk_i), .Q(reg_file[703]), .QN(
        n4388) );
  DFF_X1 reg_file_reg_9__31_ ( .D(n1809), .CK(clk_i), .Q(reg_file[735]), .QN(
        n4387) );
  DFF_X1 reg_file_reg_8__31_ ( .D(n1810), .CK(clk_i), .Q(reg_file[767]), .QN(
        n4697) );
  DFF_X1 reg_file_reg_7__31_ ( .D(n1811), .CK(clk_i), .Q(reg_file[799]), .QN(
        n4701) );
  DFF_X1 reg_file_reg_6__31_ ( .D(n1812), .CK(clk_i), .Q(reg_file[831]), .QN(
        n4177) );
  DFF_X1 reg_file_reg_5__31_ ( .D(n1813), .CK(clk_i), .Q(reg_file[863]), .QN(
        n4176) );
  DFF_X1 reg_file_reg_4__31_ ( .D(n1814), .CK(clk_i), .Q(reg_file[895]), .QN(
        n4700) );
  DFF_X1 reg_file_reg_3__31_ ( .D(n1815), .CK(clk_i), .Q(reg_file[927]), .QN(
        n4386) );
  DFF_X1 reg_file_reg_2__31_ ( .D(n1816), .CK(clk_i), .Q(reg_file[959]), .QN(
        n4385) );
  DFF_X1 reg_file_reg_1__31_ ( .D(n1817), .CK(clk_i), .Q(reg_file[991]), .QN(
        n4384) );
  DFF_X1 reg_file_reg_0__31_ ( .D(n1818), .CK(clk_i), .Q(reg_file[1023]), .QN(
        n4696) );
  DFF_X1 reg_file_reg_31__27_ ( .D(n1915), .CK(clk_i), .Q(reg_file[27]), .QN(
        n4659) );
  DFF_X1 reg_file_reg_30__27_ ( .D(n1916), .CK(clk_i), .Q(reg_file[59]), .QN(
        n4139) );
  DFF_X1 reg_file_reg_29__27_ ( .D(n1917), .CK(clk_i), .Q(reg_file[91]), .QN(
        n4138) );
  DFF_X1 reg_file_reg_28__27_ ( .D(n1918), .CK(clk_i), .Q(reg_file[123]), .QN(
        n4658) );
  DFF_X1 reg_file_reg_27__27_ ( .D(n1919), .CK(clk_i), .Q(reg_file[155]), .QN(
        n4359) );
  DFF_X1 reg_file_reg_26__27_ ( .D(n1920), .CK(clk_i), .Q(reg_file[187]), .QN(
        n4358) );
  DFF_X1 reg_file_reg_25__27_ ( .D(n1921), .CK(clk_i), .Q(reg_file[219]), .QN(
        n4657) );
  DFF_X1 reg_file_reg_24__27_ ( .D(n1922), .CK(clk_i), .Q(reg_file[251]), .QN(
        n4137) );
  DFF_X1 reg_file_reg_23__27_ ( .D(n1923), .CK(clk_i), .Q(reg_file[283]), .QN(
        n4656) );
  DFF_X1 reg_file_reg_22__27_ ( .D(n1924), .CK(clk_i), .Q(reg_file[315]), .QN(
        n4136) );
  DFF_X1 reg_file_reg_21__27_ ( .D(n1925), .CK(clk_i), .Q(reg_file[347]), .QN(
        n4135) );
  DFF_X1 reg_file_reg_20__27_ ( .D(n1926), .CK(clk_i), .Q(reg_file[379]), .QN(
        n4655) );
  DFF_X1 reg_file_reg_19__27_ ( .D(n1927), .CK(clk_i), .Q(reg_file[411]), .QN(
        n4357) );
  DFF_X1 reg_file_reg_18__27_ ( .D(n1928), .CK(clk_i), .Q(reg_file[443]), .QN(
        n4356) );
  DFF_X1 reg_file_reg_17__27_ ( .D(n1929), .CK(clk_i), .Q(reg_file[475]), .QN(
        n4654) );
  DFF_X1 reg_file_reg_16__27_ ( .D(n1930), .CK(clk_i), .Q(reg_file[507]), .QN(
        n4134) );
  DFF_X1 reg_file_reg_15__27_ ( .D(n1931), .CK(clk_i), .Q(reg_file[539]), .QN(
        n4653) );
  DFF_X1 reg_file_reg_14__27_ ( .D(n1932), .CK(clk_i), .Q(reg_file[571]), .QN(
        n4133) );
  DFF_X1 reg_file_reg_13__27_ ( .D(n1933), .CK(clk_i), .Q(reg_file[603]), .QN(
        n4132) );
  DFF_X1 reg_file_reg_12__27_ ( .D(n1934), .CK(clk_i), .Q(reg_file[635]), .QN(
        n4652) );
  DFF_X1 reg_file_reg_11__27_ ( .D(n1935), .CK(clk_i), .Q(reg_file[667]), .QN(
        n4355) );
  DFF_X1 reg_file_reg_10__27_ ( .D(n1936), .CK(clk_i), .Q(reg_file[699]), .QN(
        n4354) );
  DFF_X1 reg_file_reg_9__27_ ( .D(n1937), .CK(clk_i), .Q(reg_file[731]), .QN(
        n4651) );
  DFF_X1 reg_file_reg_8__27_ ( .D(n1938), .CK(clk_i), .Q(reg_file[763]), .QN(
        n4131) );
  DFF_X1 reg_file_reg_7__27_ ( .D(n1939), .CK(clk_i), .Q(reg_file[795]), .QN(
        n4650) );
  DFF_X1 reg_file_reg_6__27_ ( .D(n1940), .CK(clk_i), .Q(reg_file[827]), .QN(
        n4130) );
  DFF_X1 reg_file_reg_5__27_ ( .D(n1941), .CK(clk_i), .Q(reg_file[859]), .QN(
        n4129) );
  DFF_X1 reg_file_reg_4__27_ ( .D(n1942), .CK(clk_i), .Q(reg_file[891]), .QN(
        n4649) );
  DFF_X1 reg_file_reg_3__27_ ( .D(n1943), .CK(clk_i), .Q(reg_file[923]), .QN(
        n4353) );
  DFF_X1 reg_file_reg_2__27_ ( .D(n1944), .CK(clk_i), .Q(reg_file[955]), .QN(
        n4352) );
  DFF_X1 reg_file_reg_1__27_ ( .D(n1945), .CK(clk_i), .Q(reg_file[987]), .QN(
        n4648) );
  DFF_X1 reg_file_reg_0__27_ ( .D(n1946), .CK(clk_i), .Q(reg_file[1019]), .QN(
        n4128) );
  DFF_X1 reg_file_reg_31__23_ ( .D(n2043), .CK(clk_i), .Q(reg_file[23]), .QN(
        n4611) );
  DFF_X1 reg_file_reg_30__23_ ( .D(n2044), .CK(clk_i), .Q(reg_file[55]), .QN(
        n4091) );
  DFF_X1 reg_file_reg_29__23_ ( .D(n2045), .CK(clk_i), .Q(reg_file[87]), .QN(
        n4090) );
  DFF_X1 reg_file_reg_28__23_ ( .D(n2046), .CK(clk_i), .Q(reg_file[119]), .QN(
        n4610) );
  DFF_X1 reg_file_reg_27__23_ ( .D(n2047), .CK(clk_i), .Q(reg_file[151]), .QN(
        n4327) );
  DFF_X1 reg_file_reg_26__23_ ( .D(n2048), .CK(clk_i), .Q(reg_file[183]), .QN(
        n4326) );
  DFF_X1 reg_file_reg_25__23_ ( .D(n2049), .CK(clk_i), .Q(reg_file[215]), .QN(
        n4609) );
  DFF_X1 reg_file_reg_24__23_ ( .D(n2050), .CK(clk_i), .Q(reg_file[247]), .QN(
        n4089) );
  DFF_X1 reg_file_reg_23__23_ ( .D(n2051), .CK(clk_i), .Q(reg_file[279]), .QN(
        n4608) );
  DFF_X1 reg_file_reg_22__23_ ( .D(n2052), .CK(clk_i), .Q(reg_file[311]), .QN(
        n4088) );
  DFF_X1 reg_file_reg_21__23_ ( .D(n2053), .CK(clk_i), .Q(reg_file[343]), .QN(
        n4087) );
  DFF_X1 reg_file_reg_20__23_ ( .D(n2054), .CK(clk_i), .Q(reg_file[375]), .QN(
        n4607) );
  DFF_X1 reg_file_reg_19__23_ ( .D(n2055), .CK(clk_i), .Q(reg_file[407]), .QN(
        n4325) );
  DFF_X1 reg_file_reg_18__23_ ( .D(n2056), .CK(clk_i), .Q(reg_file[439]), .QN(
        n4324) );
  DFF_X1 reg_file_reg_17__23_ ( .D(n2057), .CK(clk_i), .Q(reg_file[471]), .QN(
        n4606) );
  DFF_X1 reg_file_reg_16__23_ ( .D(n2058), .CK(clk_i), .Q(reg_file[503]), .QN(
        n4086) );
  DFF_X1 reg_file_reg_15__23_ ( .D(n2059), .CK(clk_i), .Q(reg_file[535]), .QN(
        n4605) );
  DFF_X1 reg_file_reg_14__23_ ( .D(n2060), .CK(clk_i), .Q(reg_file[567]), .QN(
        n4085) );
  DFF_X1 reg_file_reg_13__23_ ( .D(n2061), .CK(clk_i), .Q(reg_file[599]), .QN(
        n4084) );
  DFF_X1 reg_file_reg_12__23_ ( .D(n2062), .CK(clk_i), .Q(reg_file[631]), .QN(
        n4604) );
  DFF_X1 reg_file_reg_11__23_ ( .D(n2063), .CK(clk_i), .Q(reg_file[663]), .QN(
        n4323) );
  DFF_X1 reg_file_reg_10__23_ ( .D(n2064), .CK(clk_i), .Q(reg_file[695]), .QN(
        n4322) );
  DFF_X1 reg_file_reg_9__23_ ( .D(n2065), .CK(clk_i), .Q(reg_file[727]), .QN(
        n4603) );
  DFF_X1 reg_file_reg_8__23_ ( .D(n2066), .CK(clk_i), .Q(reg_file[759]), .QN(
        n4083) );
  DFF_X1 reg_file_reg_7__23_ ( .D(n2067), .CK(clk_i), .Q(reg_file[791]), .QN(
        n4602) );
  DFF_X1 reg_file_reg_6__23_ ( .D(n2068), .CK(clk_i), .Q(reg_file[823]), .QN(
        n4082) );
  DFF_X1 reg_file_reg_5__23_ ( .D(n2069), .CK(clk_i), .Q(reg_file[855]), .QN(
        n4081) );
  DFF_X1 reg_file_reg_4__23_ ( .D(n2070), .CK(clk_i), .Q(reg_file[887]), .QN(
        n4601) );
  DFF_X1 reg_file_reg_3__23_ ( .D(n2071), .CK(clk_i), .Q(reg_file[919]), .QN(
        n4321) );
  DFF_X1 reg_file_reg_2__23_ ( .D(n2072), .CK(clk_i), .Q(reg_file[951]), .QN(
        n4320) );
  DFF_X1 reg_file_reg_1__23_ ( .D(n2073), .CK(clk_i), .Q(reg_file[983]), .QN(
        n4600) );
  DFF_X1 reg_file_reg_0__23_ ( .D(n2074), .CK(clk_i), .Q(reg_file[1015]), .QN(
        n4080) );
  DFF_X1 reg_file_reg_31__19_ ( .D(n2171), .CK(clk_i), .Q(reg_file[19]), .QN(
        n4563) );
  DFF_X1 reg_file_reg_30__19_ ( .D(n2172), .CK(clk_i), .Q(reg_file[51]), .QN(
        n4043) );
  DFF_X1 reg_file_reg_29__19_ ( .D(n2173), .CK(clk_i), .Q(reg_file[83]), .QN(
        n4042) );
  DFF_X1 reg_file_reg_28__19_ ( .D(n2174), .CK(clk_i), .Q(reg_file[115]), .QN(
        n4562) );
  DFF_X1 reg_file_reg_27__19_ ( .D(n2175), .CK(clk_i), .Q(reg_file[147]), .QN(
        n4295) );
  DFF_X1 reg_file_reg_26__19_ ( .D(n2176), .CK(clk_i), .Q(reg_file[179]), .QN(
        n4294) );
  DFF_X1 reg_file_reg_25__19_ ( .D(n2177), .CK(clk_i), .Q(reg_file[211]), .QN(
        n4561) );
  DFF_X1 reg_file_reg_24__19_ ( .D(n2178), .CK(clk_i), .Q(reg_file[243]), .QN(
        n4041) );
  DFF_X1 reg_file_reg_23__19_ ( .D(n2179), .CK(clk_i), .Q(reg_file[275]), .QN(
        n4560) );
  DFF_X1 reg_file_reg_22__19_ ( .D(n2180), .CK(clk_i), .Q(reg_file[307]), .QN(
        n4040) );
  DFF_X1 reg_file_reg_21__19_ ( .D(n2181), .CK(clk_i), .Q(reg_file[339]), .QN(
        n4039) );
  DFF_X1 reg_file_reg_20__19_ ( .D(n2182), .CK(clk_i), .Q(reg_file[371]), .QN(
        n4559) );
  DFF_X1 reg_file_reg_19__19_ ( .D(n2183), .CK(clk_i), .Q(reg_file[403]), .QN(
        n4293) );
  DFF_X1 reg_file_reg_18__19_ ( .D(n2184), .CK(clk_i), .Q(reg_file[435]), .QN(
        n4292) );
  DFF_X1 reg_file_reg_17__19_ ( .D(n2185), .CK(clk_i), .Q(reg_file[467]), .QN(
        n4558) );
  DFF_X1 reg_file_reg_16__19_ ( .D(n2186), .CK(clk_i), .Q(reg_file[499]), .QN(
        n4038) );
  DFF_X1 reg_file_reg_15__19_ ( .D(n2187), .CK(clk_i), .Q(reg_file[531]), .QN(
        n4557) );
  DFF_X1 reg_file_reg_14__19_ ( .D(n2188), .CK(clk_i), .Q(reg_file[563]), .QN(
        n4037) );
  DFF_X1 reg_file_reg_13__19_ ( .D(n2189), .CK(clk_i), .Q(reg_file[595]), .QN(
        n4036) );
  DFF_X1 reg_file_reg_12__19_ ( .D(n2190), .CK(clk_i), .Q(reg_file[627]), .QN(
        n4556) );
  DFF_X1 reg_file_reg_11__19_ ( .D(n2191), .CK(clk_i), .Q(reg_file[659]), .QN(
        n4291) );
  DFF_X1 reg_file_reg_10__19_ ( .D(n2192), .CK(clk_i), .Q(reg_file[691]), .QN(
        n4290) );
  DFF_X1 reg_file_reg_9__19_ ( .D(n2193), .CK(clk_i), .Q(reg_file[723]), .QN(
        n4555) );
  DFF_X1 reg_file_reg_8__19_ ( .D(n2194), .CK(clk_i), .Q(reg_file[755]), .QN(
        n4035) );
  DFF_X1 reg_file_reg_7__19_ ( .D(n2195), .CK(clk_i), .Q(reg_file[787]), .QN(
        n4554) );
  DFF_X1 reg_file_reg_6__19_ ( .D(n2196), .CK(clk_i), .Q(reg_file[819]), .QN(
        n4034) );
  DFF_X1 reg_file_reg_5__19_ ( .D(n2197), .CK(clk_i), .Q(reg_file[851]), .QN(
        n4033) );
  DFF_X1 reg_file_reg_4__19_ ( .D(n2198), .CK(clk_i), .Q(reg_file[883]), .QN(
        n4553) );
  DFF_X1 reg_file_reg_3__19_ ( .D(n2199), .CK(clk_i), .Q(reg_file[915]), .QN(
        n4289) );
  DFF_X1 reg_file_reg_2__19_ ( .D(n2200), .CK(clk_i), .Q(reg_file[947]), .QN(
        n4288) );
  DFF_X1 reg_file_reg_1__19_ ( .D(n2201), .CK(clk_i), .Q(reg_file[979]), .QN(
        n4552) );
  DFF_X1 reg_file_reg_0__19_ ( .D(n2202), .CK(clk_i), .Q(reg_file[1011]), .QN(
        n4032) );
  DFF_X1 reg_file_reg_31__13_ ( .D(n2363), .CK(clk_i), .Q(reg_file[13]), .QN(
        n4491) );
  DFF_X1 reg_file_reg_30__13_ ( .D(n2364), .CK(clk_i), .Q(reg_file[45]), .QN(
        n3971) );
  DFF_X1 reg_file_reg_29__13_ ( .D(n2365), .CK(clk_i), .Q(reg_file[77]), .QN(
        n3970) );
  DFF_X1 reg_file_reg_28__13_ ( .D(n2366), .CK(clk_i), .Q(reg_file[109]), .QN(
        n4490) );
  DFF_X1 reg_file_reg_27__13_ ( .D(n2367), .CK(clk_i), .Q(reg_file[141]), .QN(
        n4247) );
  DFF_X1 reg_file_reg_26__13_ ( .D(n2368), .CK(clk_i), .Q(reg_file[173]), .QN(
        n4246) );
  DFF_X1 reg_file_reg_25__13_ ( .D(n2369), .CK(clk_i), .Q(reg_file[205]), .QN(
        n4489) );
  DFF_X1 reg_file_reg_24__13_ ( .D(n2370), .CK(clk_i), .Q(reg_file[237]), .QN(
        n3969) );
  DFF_X1 reg_file_reg_23__13_ ( .D(n2371), .CK(clk_i), .Q(reg_file[269]), .QN(
        n4488) );
  DFF_X1 reg_file_reg_22__13_ ( .D(n2372), .CK(clk_i), .Q(reg_file[301]), .QN(
        n3968) );
  DFF_X1 reg_file_reg_21__13_ ( .D(n2373), .CK(clk_i), .Q(reg_file[333]), .QN(
        n3967) );
  DFF_X1 reg_file_reg_20__13_ ( .D(n2374), .CK(clk_i), .Q(reg_file[365]), .QN(
        n4487) );
  DFF_X1 reg_file_reg_19__13_ ( .D(n2375), .CK(clk_i), .Q(reg_file[397]), .QN(
        n4245) );
  DFF_X1 reg_file_reg_18__13_ ( .D(n2376), .CK(clk_i), .Q(reg_file[429]), .QN(
        n4244) );
  DFF_X1 reg_file_reg_17__13_ ( .D(n2377), .CK(clk_i), .Q(reg_file[461]), .QN(
        n4486) );
  DFF_X1 reg_file_reg_16__13_ ( .D(n2378), .CK(clk_i), .Q(reg_file[493]), .QN(
        n3966) );
  DFF_X1 reg_file_reg_15__13_ ( .D(n2379), .CK(clk_i), .Q(reg_file[525]), .QN(
        n4485) );
  DFF_X1 reg_file_reg_14__13_ ( .D(n2380), .CK(clk_i), .Q(reg_file[557]), .QN(
        n3965) );
  DFF_X1 reg_file_reg_13__13_ ( .D(n2381), .CK(clk_i), .Q(reg_file[589]), .QN(
        n3964) );
  DFF_X1 reg_file_reg_12__13_ ( .D(n2382), .CK(clk_i), .Q(reg_file[621]), .QN(
        n4484) );
  DFF_X1 reg_file_reg_11__13_ ( .D(n2383), .CK(clk_i), .Q(reg_file[653]), .QN(
        n4243) );
  DFF_X1 reg_file_reg_10__13_ ( .D(n2384), .CK(clk_i), .Q(reg_file[685]), .QN(
        n4242) );
  DFF_X1 reg_file_reg_9__13_ ( .D(n2385), .CK(clk_i), .Q(reg_file[717]), .QN(
        n4483) );
  DFF_X1 reg_file_reg_8__13_ ( .D(n2386), .CK(clk_i), .Q(reg_file[749]), .QN(
        n3963) );
  DFF_X1 reg_file_reg_7__13_ ( .D(n2387), .CK(clk_i), .Q(reg_file[781]), .QN(
        n4482) );
  DFF_X1 reg_file_reg_6__13_ ( .D(n2388), .CK(clk_i), .Q(reg_file[813]), .QN(
        n3962) );
  DFF_X1 reg_file_reg_5__13_ ( .D(n2389), .CK(clk_i), .Q(reg_file[845]), .QN(
        n3961) );
  DFF_X1 reg_file_reg_4__13_ ( .D(n2390), .CK(clk_i), .Q(reg_file[877]), .QN(
        n4481) );
  DFF_X1 reg_file_reg_3__13_ ( .D(n2391), .CK(clk_i), .Q(reg_file[909]), .QN(
        n4241) );
  DFF_X1 reg_file_reg_2__13_ ( .D(n2392), .CK(clk_i), .Q(reg_file[941]), .QN(
        n4240) );
  DFF_X1 reg_file_reg_1__13_ ( .D(n2393), .CK(clk_i), .Q(reg_file[973]), .QN(
        n4480) );
  DFF_X1 reg_file_reg_0__13_ ( .D(n2394), .CK(clk_i), .Q(reg_file[1005]), .QN(
        n3960) );
  DFF_X1 reg_file_reg_31__9_ ( .D(n2491), .CK(clk_i), .Q(reg_file[9]), .QN(
        n4443) );
  DFF_X1 reg_file_reg_30__9_ ( .D(n2492), .CK(clk_i), .Q(reg_file[41]), .QN(
        n3923) );
  DFF_X1 reg_file_reg_29__9_ ( .D(n2493), .CK(clk_i), .Q(reg_file[73]), .QN(
        n3922) );
  DFF_X1 reg_file_reg_28__9_ ( .D(n2494), .CK(clk_i), .Q(reg_file[105]), .QN(
        n4442) );
  DFF_X1 reg_file_reg_27__9_ ( .D(n2495), .CK(clk_i), .Q(reg_file[137]), .QN(
        n4215) );
  DFF_X1 reg_file_reg_26__9_ ( .D(n2496), .CK(clk_i), .Q(reg_file[169]), .QN(
        n4214) );
  DFF_X1 reg_file_reg_25__9_ ( .D(n2497), .CK(clk_i), .Q(reg_file[201]), .QN(
        n4441) );
  DFF_X1 reg_file_reg_24__9_ ( .D(n2498), .CK(clk_i), .Q(reg_file[233]), .QN(
        n3921) );
  DFF_X1 reg_file_reg_23__9_ ( .D(n2499), .CK(clk_i), .Q(reg_file[265]), .QN(
        n4440) );
  DFF_X1 reg_file_reg_22__9_ ( .D(n2500), .CK(clk_i), .Q(reg_file[297]), .QN(
        n3920) );
  DFF_X1 reg_file_reg_21__9_ ( .D(n2501), .CK(clk_i), .Q(reg_file[329]), .QN(
        n3919) );
  DFF_X1 reg_file_reg_20__9_ ( .D(n2502), .CK(clk_i), .Q(reg_file[361]), .QN(
        n4439) );
  DFF_X1 reg_file_reg_19__9_ ( .D(n2503), .CK(clk_i), .Q(reg_file[393]), .QN(
        n4213) );
  DFF_X1 reg_file_reg_18__9_ ( .D(n2504), .CK(clk_i), .Q(reg_file[425]), .QN(
        n4212) );
  DFF_X1 reg_file_reg_17__9_ ( .D(n2505), .CK(clk_i), .Q(reg_file[457]), .QN(
        n4438) );
  DFF_X1 reg_file_reg_16__9_ ( .D(n2506), .CK(clk_i), .Q(reg_file[489]), .QN(
        n3918) );
  DFF_X1 reg_file_reg_15__9_ ( .D(n2507), .CK(clk_i), .Q(reg_file[521]), .QN(
        n4437) );
  DFF_X1 reg_file_reg_14__9_ ( .D(n2508), .CK(clk_i), .Q(reg_file[553]), .QN(
        n3917) );
  DFF_X1 reg_file_reg_13__9_ ( .D(n2509), .CK(clk_i), .Q(reg_file[585]), .QN(
        n3916) );
  DFF_X1 reg_file_reg_12__9_ ( .D(n2510), .CK(clk_i), .Q(reg_file[617]), .QN(
        n4436) );
  DFF_X1 reg_file_reg_11__9_ ( .D(n2511), .CK(clk_i), .Q(reg_file[649]), .QN(
        n4211) );
  DFF_X1 reg_file_reg_10__9_ ( .D(n2512), .CK(clk_i), .Q(reg_file[681]), .QN(
        n4210) );
  DFF_X1 reg_file_reg_9__9_ ( .D(n2513), .CK(clk_i), .Q(reg_file[713]), .QN(
        n4435) );
  DFF_X1 reg_file_reg_8__9_ ( .D(n2514), .CK(clk_i), .Q(reg_file[745]), .QN(
        n3915) );
  DFF_X1 reg_file_reg_7__9_ ( .D(n2515), .CK(clk_i), .Q(reg_file[777]), .QN(
        n4434) );
  DFF_X1 reg_file_reg_6__9_ ( .D(n2516), .CK(clk_i), .Q(reg_file[809]), .QN(
        n3914) );
  DFF_X1 reg_file_reg_5__9_ ( .D(n2517), .CK(clk_i), .Q(reg_file[841]), .QN(
        n3913) );
  DFF_X1 reg_file_reg_4__9_ ( .D(n2518), .CK(clk_i), .Q(reg_file[873]), .QN(
        n4433) );
  DFF_X1 reg_file_reg_3__9_ ( .D(n2519), .CK(clk_i), .Q(reg_file[905]), .QN(
        n4209) );
  DFF_X1 reg_file_reg_2__9_ ( .D(n2520), .CK(clk_i), .Q(reg_file[937]), .QN(
        n4208) );
  DFF_X1 reg_file_reg_1__9_ ( .D(n2521), .CK(clk_i), .Q(reg_file[969]), .QN(
        n4432) );
  DFF_X1 reg_file_reg_0__9_ ( .D(n2522), .CK(clk_i), .Q(reg_file[1001]), .QN(
        n3912) );
  DFF_X1 reg_file_reg_31__5_ ( .D(n2619), .CK(clk_i), .Q(reg_file[5]) );
  DFF_X1 reg_file_reg_30__5_ ( .D(n2620), .CK(clk_i), .Q(reg_file[37]) );
  DFF_X1 reg_file_reg_29__5_ ( .D(n2621), .CK(clk_i), .Q(reg_file[69]) );
  DFF_X1 reg_file_reg_28__5_ ( .D(n2622), .CK(clk_i), .Q(reg_file[101]) );
  DFF_X1 reg_file_reg_27__5_ ( .D(n2623), .CK(clk_i), .Q(reg_file[133]) );
  DFF_X1 reg_file_reg_26__5_ ( .D(n2624), .CK(clk_i), .Q(reg_file[165]) );
  DFF_X1 reg_file_reg_25__5_ ( .D(n2625), .CK(clk_i), .Q(reg_file[197]) );
  DFF_X1 reg_file_reg_24__5_ ( .D(n2626), .CK(clk_i), .Q(reg_file[229]) );
  DFF_X1 reg_file_reg_23__5_ ( .D(n2627), .CK(clk_i), .Q(reg_file[261]) );
  DFF_X1 reg_file_reg_22__5_ ( .D(n2628), .CK(clk_i), .Q(reg_file[293]) );
  DFF_X1 reg_file_reg_21__5_ ( .D(n2629), .CK(clk_i), .Q(reg_file[325]) );
  DFF_X1 reg_file_reg_20__5_ ( .D(n2630), .CK(clk_i), .Q(reg_file[357]) );
  DFF_X1 reg_file_reg_19__5_ ( .D(n2631), .CK(clk_i), .Q(reg_file[389]) );
  DFF_X1 reg_file_reg_18__5_ ( .D(n2632), .CK(clk_i), .Q(reg_file[421]) );
  DFF_X1 reg_file_reg_17__5_ ( .D(n2633), .CK(clk_i), .Q(reg_file[453]) );
  DFF_X1 reg_file_reg_16__5_ ( .D(n2634), .CK(clk_i), .Q(reg_file[485]) );
  DFF_X1 reg_file_reg_15__5_ ( .D(n2635), .CK(clk_i), .Q(reg_file[517]) );
  DFF_X1 reg_file_reg_14__5_ ( .D(n2636), .CK(clk_i), .Q(reg_file[549]) );
  DFF_X1 reg_file_reg_13__5_ ( .D(n2637), .CK(clk_i), .Q(reg_file[581]) );
  DFF_X1 reg_file_reg_12__5_ ( .D(n2638), .CK(clk_i), .Q(reg_file[613]) );
  DFF_X1 reg_file_reg_11__5_ ( .D(n2639), .CK(clk_i), .Q(reg_file[645]) );
  DFF_X1 reg_file_reg_10__5_ ( .D(n2640), .CK(clk_i), .Q(reg_file[677]) );
  DFF_X1 reg_file_reg_9__5_ ( .D(n2641), .CK(clk_i), .Q(reg_file[709]) );
  DFF_X1 reg_file_reg_8__5_ ( .D(n2642), .CK(clk_i), .Q(reg_file[741]) );
  DFF_X1 reg_file_reg_7__5_ ( .D(n2643), .CK(clk_i), .Q(reg_file[773]) );
  DFF_X1 reg_file_reg_6__5_ ( .D(n2644), .CK(clk_i), .Q(reg_file[805]) );
  DFF_X1 reg_file_reg_5__5_ ( .D(n2645), .CK(clk_i), .Q(reg_file[837]) );
  DFF_X1 reg_file_reg_4__5_ ( .D(n2646), .CK(clk_i), .Q(reg_file[869]) );
  DFF_X1 reg_file_reg_3__5_ ( .D(n2647), .CK(clk_i), .Q(reg_file[901]) );
  DFF_X1 reg_file_reg_2__5_ ( .D(n2648), .CK(clk_i), .Q(reg_file[933]) );
  DFF_X1 reg_file_reg_1__5_ ( .D(n2649), .CK(clk_i), .Q(reg_file[965]) );
  DFF_X1 reg_file_reg_0__5_ ( .D(n2650), .CK(clk_i), .Q(reg_file[997]) );
  DFF_X1 reg_file_reg_31__1_ ( .D(n2747), .CK(clk_i), .Q(reg_file[1]) );
  DFF_X1 reg_file_reg_30__1_ ( .D(n2748), .CK(clk_i), .Q(reg_file[33]) );
  DFF_X1 reg_file_reg_29__1_ ( .D(n2749), .CK(clk_i), .Q(reg_file[65]) );
  DFF_X1 reg_file_reg_28__1_ ( .D(n2750), .CK(clk_i), .Q(reg_file[97]) );
  DFF_X1 reg_file_reg_27__1_ ( .D(n2751), .CK(clk_i), .Q(reg_file[129]) );
  DFF_X1 reg_file_reg_26__1_ ( .D(n2752), .CK(clk_i), .Q(reg_file[161]) );
  DFF_X1 reg_file_reg_25__1_ ( .D(n2753), .CK(clk_i), .Q(reg_file[193]) );
  DFF_X1 reg_file_reg_24__1_ ( .D(n2754), .CK(clk_i), .Q(reg_file[225]) );
  DFF_X1 reg_file_reg_23__1_ ( .D(n2755), .CK(clk_i), .Q(reg_file[257]) );
  DFF_X1 reg_file_reg_22__1_ ( .D(n2756), .CK(clk_i), .Q(reg_file[289]) );
  DFF_X1 reg_file_reg_21__1_ ( .D(n2757), .CK(clk_i), .Q(reg_file[321]) );
  DFF_X1 reg_file_reg_20__1_ ( .D(n2758), .CK(clk_i), .Q(reg_file[353]) );
  DFF_X1 reg_file_reg_19__1_ ( .D(n2759), .CK(clk_i), .Q(reg_file[385]) );
  DFF_X1 reg_file_reg_18__1_ ( .D(n2760), .CK(clk_i), .Q(reg_file[417]) );
  DFF_X1 reg_file_reg_17__1_ ( .D(n2761), .CK(clk_i), .Q(reg_file[449]) );
  DFF_X1 reg_file_reg_16__1_ ( .D(n2762), .CK(clk_i), .Q(reg_file[481]) );
  DFF_X1 reg_file_reg_15__1_ ( .D(n2763), .CK(clk_i), .Q(reg_file[513]) );
  DFF_X1 reg_file_reg_14__1_ ( .D(n2764), .CK(clk_i), .Q(reg_file[545]) );
  DFF_X1 reg_file_reg_13__1_ ( .D(n2765), .CK(clk_i), .Q(reg_file[577]) );
  DFF_X1 reg_file_reg_12__1_ ( .D(n2766), .CK(clk_i), .Q(reg_file[609]) );
  DFF_X1 reg_file_reg_11__1_ ( .D(n2767), .CK(clk_i), .Q(reg_file[641]) );
  DFF_X1 reg_file_reg_10__1_ ( .D(n2768), .CK(clk_i), .Q(reg_file[673]) );
  DFF_X1 reg_file_reg_9__1_ ( .D(n2769), .CK(clk_i), .Q(reg_file[705]) );
  DFF_X1 reg_file_reg_8__1_ ( .D(n2770), .CK(clk_i), .Q(reg_file[737]) );
  DFF_X1 reg_file_reg_7__1_ ( .D(n2771), .CK(clk_i), .Q(reg_file[769]) );
  DFF_X1 reg_file_reg_6__1_ ( .D(n2772), .CK(clk_i), .Q(reg_file[801]) );
  DFF_X1 reg_file_reg_5__1_ ( .D(n2773), .CK(clk_i), .Q(reg_file[833]) );
  DFF_X1 reg_file_reg_4__1_ ( .D(n2774), .CK(clk_i), .Q(reg_file[865]) );
  DFF_X1 reg_file_reg_3__1_ ( .D(n2775), .CK(clk_i), .Q(reg_file[897]) );
  DFF_X1 reg_file_reg_2__1_ ( .D(n2776), .CK(clk_i), .Q(reg_file[929]) );
  DFF_X1 reg_file_reg_1__1_ ( .D(n2777), .CK(clk_i), .Q(reg_file[961]) );
  DFF_X1 reg_file_reg_0__1_ ( .D(n2778), .CK(clk_i), .Q(reg_file[993]) );
  DFF_X1 reg_file_reg_31__30_ ( .D(n1819), .CK(clk_i), .Q(reg_file[30]), .QN(
        n4695) );
  DFF_X1 reg_file_reg_30__30_ ( .D(n1820), .CK(clk_i), .Q(reg_file[62]), .QN(
        n4175) );
  DFF_X1 reg_file_reg_29__30_ ( .D(n1821), .CK(clk_i), .Q(reg_file[94]), .QN(
        n4174) );
  DFF_X1 reg_file_reg_28__30_ ( .D(n1822), .CK(clk_i), .Q(reg_file[126]), .QN(
        n4694) );
  DFF_X1 reg_file_reg_27__30_ ( .D(n1823), .CK(clk_i), .Q(reg_file[158]), .QN(
        n4383) );
  DFF_X1 reg_file_reg_26__30_ ( .D(n1824), .CK(clk_i), .Q(reg_file[190]), .QN(
        n4382) );
  DFF_X1 reg_file_reg_25__30_ ( .D(n1825), .CK(clk_i), .Q(reg_file[222]), .QN(
        n4693) );
  DFF_X1 reg_file_reg_24__30_ ( .D(n1826), .CK(clk_i), .Q(reg_file[254]), .QN(
        n4173) );
  DFF_X1 reg_file_reg_23__30_ ( .D(n1827), .CK(clk_i), .Q(reg_file[286]), .QN(
        n4692) );
  DFF_X1 reg_file_reg_22__30_ ( .D(n1828), .CK(clk_i), .Q(reg_file[318]), .QN(
        n4172) );
  DFF_X1 reg_file_reg_21__30_ ( .D(n1829), .CK(clk_i), .Q(reg_file[350]), .QN(
        n4171) );
  DFF_X1 reg_file_reg_20__30_ ( .D(n1830), .CK(clk_i), .Q(reg_file[382]), .QN(
        n4691) );
  DFF_X1 reg_file_reg_19__30_ ( .D(n1831), .CK(clk_i), .Q(reg_file[414]), .QN(
        n4381) );
  DFF_X1 reg_file_reg_18__30_ ( .D(n1832), .CK(clk_i), .Q(reg_file[446]), .QN(
        n4380) );
  DFF_X1 reg_file_reg_17__30_ ( .D(n1833), .CK(clk_i), .Q(reg_file[478]), .QN(
        n4690) );
  DFF_X1 reg_file_reg_16__30_ ( .D(n1834), .CK(clk_i), .Q(reg_file[510]), .QN(
        n4170) );
  DFF_X1 reg_file_reg_15__30_ ( .D(n1835), .CK(clk_i), .Q(reg_file[542]), .QN(
        n4689) );
  DFF_X1 reg_file_reg_14__30_ ( .D(n1836), .CK(clk_i), .Q(reg_file[574]), .QN(
        n4169) );
  DFF_X1 reg_file_reg_13__30_ ( .D(n1837), .CK(clk_i), .Q(reg_file[606]), .QN(
        n4168) );
  DFF_X1 reg_file_reg_12__30_ ( .D(n1838), .CK(clk_i), .Q(reg_file[638]), .QN(
        n4688) );
  DFF_X1 reg_file_reg_11__30_ ( .D(n1839), .CK(clk_i), .Q(reg_file[670]), .QN(
        n4379) );
  DFF_X1 reg_file_reg_10__30_ ( .D(n1840), .CK(clk_i), .Q(reg_file[702]), .QN(
        n4378) );
  DFF_X1 reg_file_reg_9__30_ ( .D(n1841), .CK(clk_i), .Q(reg_file[734]), .QN(
        n4687) );
  DFF_X1 reg_file_reg_8__30_ ( .D(n1842), .CK(clk_i), .Q(reg_file[766]), .QN(
        n4167) );
  DFF_X1 reg_file_reg_7__30_ ( .D(n1843), .CK(clk_i), .Q(reg_file[798]), .QN(
        n4686) );
  DFF_X1 reg_file_reg_6__30_ ( .D(n1844), .CK(clk_i), .Q(reg_file[830]), .QN(
        n4166) );
  DFF_X1 reg_file_reg_5__30_ ( .D(n1845), .CK(clk_i), .Q(reg_file[862]), .QN(
        n4165) );
  DFF_X1 reg_file_reg_4__30_ ( .D(n1846), .CK(clk_i), .Q(reg_file[894]), .QN(
        n4685) );
  DFF_X1 reg_file_reg_3__30_ ( .D(n1847), .CK(clk_i), .Q(reg_file[926]), .QN(
        n4377) );
  DFF_X1 reg_file_reg_2__30_ ( .D(n1848), .CK(clk_i), .Q(reg_file[958]), .QN(
        n4376) );
  DFF_X1 reg_file_reg_1__30_ ( .D(n1849), .CK(clk_i), .Q(reg_file[990]), .QN(
        n4684) );
  DFF_X1 reg_file_reg_0__30_ ( .D(n1850), .CK(clk_i), .Q(reg_file[1022]), .QN(
        n4164) );
  DFF_X1 reg_file_reg_31__26_ ( .D(n1947), .CK(clk_i), .Q(reg_file[26]), .QN(
        n4647) );
  DFF_X1 reg_file_reg_30__26_ ( .D(n1948), .CK(clk_i), .Q(reg_file[58]), .QN(
        n4127) );
  DFF_X1 reg_file_reg_29__26_ ( .D(n1949), .CK(clk_i), .Q(reg_file[90]), .QN(
        n4126) );
  DFF_X1 reg_file_reg_28__26_ ( .D(n1950), .CK(clk_i), .Q(reg_file[122]), .QN(
        n4646) );
  DFF_X1 reg_file_reg_27__26_ ( .D(n1951), .CK(clk_i), .Q(reg_file[154]), .QN(
        n4351) );
  DFF_X1 reg_file_reg_26__26_ ( .D(n1952), .CK(clk_i), .Q(reg_file[186]), .QN(
        n4350) );
  DFF_X1 reg_file_reg_25__26_ ( .D(n1953), .CK(clk_i), .Q(reg_file[218]), .QN(
        n4645) );
  DFF_X1 reg_file_reg_24__26_ ( .D(n1954), .CK(clk_i), .Q(reg_file[250]), .QN(
        n4125) );
  DFF_X1 reg_file_reg_23__26_ ( .D(n1955), .CK(clk_i), .Q(reg_file[282]), .QN(
        n4644) );
  DFF_X1 reg_file_reg_22__26_ ( .D(n1956), .CK(clk_i), .Q(reg_file[314]), .QN(
        n4124) );
  DFF_X1 reg_file_reg_21__26_ ( .D(n1957), .CK(clk_i), .Q(reg_file[346]), .QN(
        n4123) );
  DFF_X1 reg_file_reg_20__26_ ( .D(n1958), .CK(clk_i), .Q(reg_file[378]), .QN(
        n4643) );
  DFF_X1 reg_file_reg_19__26_ ( .D(n1959), .CK(clk_i), .Q(reg_file[410]), .QN(
        n4349) );
  DFF_X1 reg_file_reg_18__26_ ( .D(n1960), .CK(clk_i), .Q(reg_file[442]), .QN(
        n4348) );
  DFF_X1 reg_file_reg_17__26_ ( .D(n1961), .CK(clk_i), .Q(reg_file[474]), .QN(
        n4642) );
  DFF_X1 reg_file_reg_16__26_ ( .D(n1962), .CK(clk_i), .Q(reg_file[506]), .QN(
        n4122) );
  DFF_X1 reg_file_reg_15__26_ ( .D(n1963), .CK(clk_i), .Q(reg_file[538]), .QN(
        n4641) );
  DFF_X1 reg_file_reg_14__26_ ( .D(n1964), .CK(clk_i), .Q(reg_file[570]), .QN(
        n4121) );
  DFF_X1 reg_file_reg_13__26_ ( .D(n1965), .CK(clk_i), .Q(reg_file[602]), .QN(
        n4120) );
  DFF_X1 reg_file_reg_12__26_ ( .D(n1966), .CK(clk_i), .Q(reg_file[634]), .QN(
        n4640) );
  DFF_X1 reg_file_reg_11__26_ ( .D(n1967), .CK(clk_i), .Q(reg_file[666]), .QN(
        n4347) );
  DFF_X1 reg_file_reg_10__26_ ( .D(n1968), .CK(clk_i), .Q(reg_file[698]), .QN(
        n4346) );
  DFF_X1 reg_file_reg_9__26_ ( .D(n1969), .CK(clk_i), .Q(reg_file[730]), .QN(
        n4639) );
  DFF_X1 reg_file_reg_8__26_ ( .D(n1970), .CK(clk_i), .Q(reg_file[762]), .QN(
        n4119) );
  DFF_X1 reg_file_reg_7__26_ ( .D(n1971), .CK(clk_i), .Q(reg_file[794]), .QN(
        n4638) );
  DFF_X1 reg_file_reg_6__26_ ( .D(n1972), .CK(clk_i), .Q(reg_file[826]), .QN(
        n4118) );
  DFF_X1 reg_file_reg_5__26_ ( .D(n1973), .CK(clk_i), .Q(reg_file[858]), .QN(
        n4117) );
  DFF_X1 reg_file_reg_4__26_ ( .D(n1974), .CK(clk_i), .Q(reg_file[890]), .QN(
        n4637) );
  DFF_X1 reg_file_reg_3__26_ ( .D(n1975), .CK(clk_i), .Q(reg_file[922]), .QN(
        n4345) );
  DFF_X1 reg_file_reg_2__26_ ( .D(n1976), .CK(clk_i), .Q(reg_file[954]), .QN(
        n4344) );
  DFF_X1 reg_file_reg_1__26_ ( .D(n1977), .CK(clk_i), .Q(reg_file[986]), .QN(
        n4636) );
  DFF_X1 reg_file_reg_0__26_ ( .D(n1978), .CK(clk_i), .Q(reg_file[1018]), .QN(
        n4116) );
  DFF_X1 reg_file_reg_31__22_ ( .D(n2075), .CK(clk_i), .Q(reg_file[22]), .QN(
        n4599) );
  DFF_X1 reg_file_reg_30__22_ ( .D(n2076), .CK(clk_i), .Q(reg_file[54]), .QN(
        n4079) );
  DFF_X1 reg_file_reg_29__22_ ( .D(n2077), .CK(clk_i), .Q(reg_file[86]), .QN(
        n4078) );
  DFF_X1 reg_file_reg_28__22_ ( .D(n2078), .CK(clk_i), .Q(reg_file[118]), .QN(
        n4598) );
  DFF_X1 reg_file_reg_27__22_ ( .D(n2079), .CK(clk_i), .Q(reg_file[150]), .QN(
        n4319) );
  DFF_X1 reg_file_reg_26__22_ ( .D(n2080), .CK(clk_i), .Q(reg_file[182]), .QN(
        n4318) );
  DFF_X1 reg_file_reg_25__22_ ( .D(n2081), .CK(clk_i), .Q(reg_file[214]), .QN(
        n4597) );
  DFF_X1 reg_file_reg_24__22_ ( .D(n2082), .CK(clk_i), .Q(reg_file[246]), .QN(
        n4077) );
  DFF_X1 reg_file_reg_23__22_ ( .D(n2083), .CK(clk_i), .Q(reg_file[278]), .QN(
        n4596) );
  DFF_X1 reg_file_reg_22__22_ ( .D(n2084), .CK(clk_i), .Q(reg_file[310]), .QN(
        n4076) );
  DFF_X1 reg_file_reg_21__22_ ( .D(n2085), .CK(clk_i), .Q(reg_file[342]), .QN(
        n4075) );
  DFF_X1 reg_file_reg_20__22_ ( .D(n2086), .CK(clk_i), .Q(reg_file[374]), .QN(
        n4595) );
  DFF_X1 reg_file_reg_19__22_ ( .D(n2087), .CK(clk_i), .Q(reg_file[406]), .QN(
        n4317) );
  DFF_X1 reg_file_reg_18__22_ ( .D(n2088), .CK(clk_i), .Q(reg_file[438]), .QN(
        n4316) );
  DFF_X1 reg_file_reg_17__22_ ( .D(n2089), .CK(clk_i), .Q(reg_file[470]), .QN(
        n4594) );
  DFF_X1 reg_file_reg_16__22_ ( .D(n2090), .CK(clk_i), .Q(reg_file[502]), .QN(
        n4074) );
  DFF_X1 reg_file_reg_15__22_ ( .D(n2091), .CK(clk_i), .Q(reg_file[534]), .QN(
        n4593) );
  DFF_X1 reg_file_reg_14__22_ ( .D(n2092), .CK(clk_i), .Q(reg_file[566]), .QN(
        n4073) );
  DFF_X1 reg_file_reg_13__22_ ( .D(n2093), .CK(clk_i), .Q(reg_file[598]), .QN(
        n4072) );
  DFF_X1 reg_file_reg_12__22_ ( .D(n2094), .CK(clk_i), .Q(reg_file[630]), .QN(
        n4592) );
  DFF_X1 reg_file_reg_11__22_ ( .D(n2095), .CK(clk_i), .Q(reg_file[662]), .QN(
        n4315) );
  DFF_X1 reg_file_reg_10__22_ ( .D(n2096), .CK(clk_i), .Q(reg_file[694]), .QN(
        n4314) );
  DFF_X1 reg_file_reg_9__22_ ( .D(n2097), .CK(clk_i), .Q(reg_file[726]), .QN(
        n4591) );
  DFF_X1 reg_file_reg_8__22_ ( .D(n2098), .CK(clk_i), .Q(reg_file[758]), .QN(
        n4071) );
  DFF_X1 reg_file_reg_7__22_ ( .D(n2099), .CK(clk_i), .Q(reg_file[790]), .QN(
        n4590) );
  DFF_X1 reg_file_reg_6__22_ ( .D(n2100), .CK(clk_i), .Q(reg_file[822]), .QN(
        n4070) );
  DFF_X1 reg_file_reg_5__22_ ( .D(n2101), .CK(clk_i), .Q(reg_file[854]), .QN(
        n4069) );
  DFF_X1 reg_file_reg_4__22_ ( .D(n2102), .CK(clk_i), .Q(reg_file[886]), .QN(
        n4589) );
  DFF_X1 reg_file_reg_3__22_ ( .D(n2103), .CK(clk_i), .Q(reg_file[918]), .QN(
        n4313) );
  DFF_X1 reg_file_reg_2__22_ ( .D(n2104), .CK(clk_i), .Q(reg_file[950]), .QN(
        n4312) );
  DFF_X1 reg_file_reg_1__22_ ( .D(n2105), .CK(clk_i), .Q(reg_file[982]), .QN(
        n4588) );
  DFF_X1 reg_file_reg_0__22_ ( .D(n2106), .CK(clk_i), .Q(reg_file[1014]), .QN(
        n4068) );
  DFF_X1 reg_file_reg_31__18_ ( .D(n2203), .CK(clk_i), .Q(reg_file[18]), .QN(
        n4551) );
  DFF_X1 reg_file_reg_30__18_ ( .D(n2204), .CK(clk_i), .Q(reg_file[50]), .QN(
        n4031) );
  DFF_X1 reg_file_reg_29__18_ ( .D(n2205), .CK(clk_i), .Q(reg_file[82]), .QN(
        n4030) );
  DFF_X1 reg_file_reg_28__18_ ( .D(n2206), .CK(clk_i), .Q(reg_file[114]), .QN(
        n4550) );
  DFF_X1 reg_file_reg_27__18_ ( .D(n2207), .CK(clk_i), .Q(reg_file[146]), .QN(
        n4287) );
  DFF_X1 reg_file_reg_26__18_ ( .D(n2208), .CK(clk_i), .Q(reg_file[178]), .QN(
        n4286) );
  DFF_X1 reg_file_reg_25__18_ ( .D(n2209), .CK(clk_i), .Q(reg_file[210]), .QN(
        n4549) );
  DFF_X1 reg_file_reg_24__18_ ( .D(n2210), .CK(clk_i), .Q(reg_file[242]), .QN(
        n4029) );
  DFF_X1 reg_file_reg_23__18_ ( .D(n2211), .CK(clk_i), .Q(reg_file[274]), .QN(
        n4548) );
  DFF_X1 reg_file_reg_22__18_ ( .D(n2212), .CK(clk_i), .Q(reg_file[306]), .QN(
        n4028) );
  DFF_X1 reg_file_reg_21__18_ ( .D(n2213), .CK(clk_i), .Q(reg_file[338]), .QN(
        n4027) );
  DFF_X1 reg_file_reg_20__18_ ( .D(n2214), .CK(clk_i), .Q(reg_file[370]), .QN(
        n4547) );
  DFF_X1 reg_file_reg_19__18_ ( .D(n2215), .CK(clk_i), .Q(reg_file[402]), .QN(
        n4285) );
  DFF_X1 reg_file_reg_18__18_ ( .D(n2216), .CK(clk_i), .Q(reg_file[434]), .QN(
        n4284) );
  DFF_X1 reg_file_reg_17__18_ ( .D(n2217), .CK(clk_i), .Q(reg_file[466]), .QN(
        n4546) );
  DFF_X1 reg_file_reg_16__18_ ( .D(n2218), .CK(clk_i), .Q(reg_file[498]), .QN(
        n4026) );
  DFF_X1 reg_file_reg_15__18_ ( .D(n2219), .CK(clk_i), .Q(reg_file[530]), .QN(
        n4545) );
  DFF_X1 reg_file_reg_14__18_ ( .D(n2220), .CK(clk_i), .Q(reg_file[562]), .QN(
        n4025) );
  DFF_X1 reg_file_reg_13__18_ ( .D(n2221), .CK(clk_i), .Q(reg_file[594]), .QN(
        n4024) );
  DFF_X1 reg_file_reg_12__18_ ( .D(n2222), .CK(clk_i), .Q(reg_file[626]), .QN(
        n4544) );
  DFF_X1 reg_file_reg_11__18_ ( .D(n2223), .CK(clk_i), .Q(reg_file[658]), .QN(
        n4283) );
  DFF_X1 reg_file_reg_10__18_ ( .D(n2224), .CK(clk_i), .Q(reg_file[690]), .QN(
        n4282) );
  DFF_X1 reg_file_reg_9__18_ ( .D(n2225), .CK(clk_i), .Q(reg_file[722]), .QN(
        n4543) );
  DFF_X1 reg_file_reg_8__18_ ( .D(n2226), .CK(clk_i), .Q(reg_file[754]), .QN(
        n4023) );
  DFF_X1 reg_file_reg_7__18_ ( .D(n2227), .CK(clk_i), .Q(reg_file[786]), .QN(
        n4542) );
  DFF_X1 reg_file_reg_6__18_ ( .D(n2228), .CK(clk_i), .Q(reg_file[818]), .QN(
        n4022) );
  DFF_X1 reg_file_reg_5__18_ ( .D(n2229), .CK(clk_i), .Q(reg_file[850]), .QN(
        n4021) );
  DFF_X1 reg_file_reg_4__18_ ( .D(n2230), .CK(clk_i), .Q(reg_file[882]), .QN(
        n4541) );
  DFF_X1 reg_file_reg_3__18_ ( .D(n2231), .CK(clk_i), .Q(reg_file[914]), .QN(
        n4281) );
  DFF_X1 reg_file_reg_2__18_ ( .D(n2232), .CK(clk_i), .Q(reg_file[946]), .QN(
        n4280) );
  DFF_X1 reg_file_reg_1__18_ ( .D(n2233), .CK(clk_i), .Q(reg_file[978]), .QN(
        n4540) );
  DFF_X1 reg_file_reg_0__18_ ( .D(n2234), .CK(clk_i), .Q(reg_file[1010]), .QN(
        n4020) );
  DFF_X1 reg_file_reg_31__14_ ( .D(n2331), .CK(clk_i), .Q(reg_file[14]), .QN(
        n4503) );
  DFF_X1 reg_file_reg_30__14_ ( .D(n2332), .CK(clk_i), .Q(reg_file[46]), .QN(
        n3983) );
  DFF_X1 reg_file_reg_29__14_ ( .D(n2333), .CK(clk_i), .Q(reg_file[78]), .QN(
        n3982) );
  DFF_X1 reg_file_reg_28__14_ ( .D(n2334), .CK(clk_i), .Q(reg_file[110]), .QN(
        n4502) );
  DFF_X1 reg_file_reg_27__14_ ( .D(n2335), .CK(clk_i), .Q(reg_file[142]), .QN(
        n4255) );
  DFF_X1 reg_file_reg_26__14_ ( .D(n2336), .CK(clk_i), .Q(reg_file[174]), .QN(
        n4254) );
  DFF_X1 reg_file_reg_25__14_ ( .D(n2337), .CK(clk_i), .Q(reg_file[206]), .QN(
        n4501) );
  DFF_X1 reg_file_reg_24__14_ ( .D(n2338), .CK(clk_i), .Q(reg_file[238]), .QN(
        n3981) );
  DFF_X1 reg_file_reg_23__14_ ( .D(n2339), .CK(clk_i), .Q(reg_file[270]), .QN(
        n4500) );
  DFF_X1 reg_file_reg_22__14_ ( .D(n2340), .CK(clk_i), .Q(reg_file[302]), .QN(
        n3980) );
  DFF_X1 reg_file_reg_21__14_ ( .D(n2341), .CK(clk_i), .Q(reg_file[334]), .QN(
        n3979) );
  DFF_X1 reg_file_reg_20__14_ ( .D(n2342), .CK(clk_i), .Q(reg_file[366]), .QN(
        n4499) );
  DFF_X1 reg_file_reg_19__14_ ( .D(n2343), .CK(clk_i), .Q(reg_file[398]), .QN(
        n4253) );
  DFF_X1 reg_file_reg_18__14_ ( .D(n2344), .CK(clk_i), .Q(reg_file[430]), .QN(
        n4252) );
  DFF_X1 reg_file_reg_17__14_ ( .D(n2345), .CK(clk_i), .Q(reg_file[462]), .QN(
        n4498) );
  DFF_X1 reg_file_reg_16__14_ ( .D(n2346), .CK(clk_i), .Q(reg_file[494]), .QN(
        n3978) );
  DFF_X1 reg_file_reg_15__14_ ( .D(n2347), .CK(clk_i), .Q(reg_file[526]), .QN(
        n4497) );
  DFF_X1 reg_file_reg_14__14_ ( .D(n2348), .CK(clk_i), .Q(reg_file[558]), .QN(
        n3977) );
  DFF_X1 reg_file_reg_13__14_ ( .D(n2349), .CK(clk_i), .Q(reg_file[590]), .QN(
        n3976) );
  DFF_X1 reg_file_reg_12__14_ ( .D(n2350), .CK(clk_i), .Q(reg_file[622]), .QN(
        n4496) );
  DFF_X1 reg_file_reg_11__14_ ( .D(n2351), .CK(clk_i), .Q(reg_file[654]), .QN(
        n4251) );
  DFF_X1 reg_file_reg_10__14_ ( .D(n2352), .CK(clk_i), .Q(reg_file[686]), .QN(
        n4250) );
  DFF_X1 reg_file_reg_9__14_ ( .D(n2353), .CK(clk_i), .Q(reg_file[718]), .QN(
        n4495) );
  DFF_X1 reg_file_reg_8__14_ ( .D(n2354), .CK(clk_i), .Q(reg_file[750]), .QN(
        n3975) );
  DFF_X1 reg_file_reg_7__14_ ( .D(n2355), .CK(clk_i), .Q(reg_file[782]), .QN(
        n4494) );
  DFF_X1 reg_file_reg_6__14_ ( .D(n2356), .CK(clk_i), .Q(reg_file[814]), .QN(
        n3974) );
  DFF_X1 reg_file_reg_5__14_ ( .D(n2357), .CK(clk_i), .Q(reg_file[846]), .QN(
        n3973) );
  DFF_X1 reg_file_reg_4__14_ ( .D(n2358), .CK(clk_i), .Q(reg_file[878]), .QN(
        n4493) );
  DFF_X1 reg_file_reg_3__14_ ( .D(n2359), .CK(clk_i), .Q(reg_file[910]), .QN(
        n4249) );
  DFF_X1 reg_file_reg_2__14_ ( .D(n2360), .CK(clk_i), .Q(reg_file[942]), .QN(
        n4248) );
  DFF_X1 reg_file_reg_1__14_ ( .D(n2361), .CK(clk_i), .Q(reg_file[974]), .QN(
        n4492) );
  DFF_X1 reg_file_reg_0__14_ ( .D(n2362), .CK(clk_i), .Q(reg_file[1006]), .QN(
        n3972) );
  DFF_X1 reg_file_reg_31__10_ ( .D(n2459), .CK(clk_i), .Q(reg_file[10]), .QN(
        n4455) );
  DFF_X1 reg_file_reg_30__10_ ( .D(n2460), .CK(clk_i), .Q(reg_file[42]), .QN(
        n3935) );
  DFF_X1 reg_file_reg_29__10_ ( .D(n2461), .CK(clk_i), .Q(reg_file[74]), .QN(
        n3934) );
  DFF_X1 reg_file_reg_28__10_ ( .D(n2462), .CK(clk_i), .Q(reg_file[106]), .QN(
        n4454) );
  DFF_X1 reg_file_reg_27__10_ ( .D(n2463), .CK(clk_i), .Q(reg_file[138]), .QN(
        n4223) );
  DFF_X1 reg_file_reg_26__10_ ( .D(n2464), .CK(clk_i), .Q(reg_file[170]), .QN(
        n4222) );
  DFF_X1 reg_file_reg_25__10_ ( .D(n2465), .CK(clk_i), .Q(reg_file[202]), .QN(
        n4453) );
  DFF_X1 reg_file_reg_24__10_ ( .D(n2466), .CK(clk_i), .Q(reg_file[234]), .QN(
        n3933) );
  DFF_X1 reg_file_reg_23__10_ ( .D(n2467), .CK(clk_i), .Q(reg_file[266]), .QN(
        n4452) );
  DFF_X1 reg_file_reg_22__10_ ( .D(n2468), .CK(clk_i), .Q(reg_file[298]), .QN(
        n3932) );
  DFF_X1 reg_file_reg_21__10_ ( .D(n2469), .CK(clk_i), .Q(reg_file[330]), .QN(
        n3931) );
  DFF_X1 reg_file_reg_20__10_ ( .D(n2470), .CK(clk_i), .Q(reg_file[362]), .QN(
        n4451) );
  DFF_X1 reg_file_reg_19__10_ ( .D(n2471), .CK(clk_i), .Q(reg_file[394]), .QN(
        n4221) );
  DFF_X1 reg_file_reg_18__10_ ( .D(n2472), .CK(clk_i), .Q(reg_file[426]), .QN(
        n4220) );
  DFF_X1 reg_file_reg_17__10_ ( .D(n2473), .CK(clk_i), .Q(reg_file[458]), .QN(
        n4450) );
  DFF_X1 reg_file_reg_16__10_ ( .D(n2474), .CK(clk_i), .Q(reg_file[490]), .QN(
        n3930) );
  DFF_X1 reg_file_reg_15__10_ ( .D(n2475), .CK(clk_i), .Q(reg_file[522]), .QN(
        n4449) );
  DFF_X1 reg_file_reg_14__10_ ( .D(n2476), .CK(clk_i), .Q(reg_file[554]), .QN(
        n3929) );
  DFF_X1 reg_file_reg_13__10_ ( .D(n2477), .CK(clk_i), .Q(reg_file[586]), .QN(
        n3928) );
  DFF_X1 reg_file_reg_12__10_ ( .D(n2478), .CK(clk_i), .Q(reg_file[618]), .QN(
        n4448) );
  DFF_X1 reg_file_reg_11__10_ ( .D(n2479), .CK(clk_i), .Q(reg_file[650]), .QN(
        n4219) );
  DFF_X1 reg_file_reg_10__10_ ( .D(n2480), .CK(clk_i), .Q(reg_file[682]), .QN(
        n4218) );
  DFF_X1 reg_file_reg_9__10_ ( .D(n2481), .CK(clk_i), .Q(reg_file[714]), .QN(
        n4447) );
  DFF_X1 reg_file_reg_8__10_ ( .D(n2482), .CK(clk_i), .Q(reg_file[746]), .QN(
        n3927) );
  DFF_X1 reg_file_reg_7__10_ ( .D(n2483), .CK(clk_i), .Q(reg_file[778]), .QN(
        n4446) );
  DFF_X1 reg_file_reg_6__10_ ( .D(n2484), .CK(clk_i), .Q(reg_file[810]), .QN(
        n3926) );
  DFF_X1 reg_file_reg_5__10_ ( .D(n2485), .CK(clk_i), .Q(reg_file[842]), .QN(
        n3925) );
  DFF_X1 reg_file_reg_4__10_ ( .D(n2486), .CK(clk_i), .Q(reg_file[874]), .QN(
        n4445) );
  DFF_X1 reg_file_reg_3__10_ ( .D(n2487), .CK(clk_i), .Q(reg_file[906]), .QN(
        n4217) );
  DFF_X1 reg_file_reg_2__10_ ( .D(n2488), .CK(clk_i), .Q(reg_file[938]), .QN(
        n4216) );
  DFF_X1 reg_file_reg_1__10_ ( .D(n2489), .CK(clk_i), .Q(reg_file[970]), .QN(
        n4444) );
  DFF_X1 reg_file_reg_0__10_ ( .D(n2490), .CK(clk_i), .Q(reg_file[1002]), .QN(
        n3924) );
  DFF_X1 reg_file_reg_31__6_ ( .D(n2587), .CK(clk_i), .Q(reg_file[6]), .QN(
        n4407) );
  DFF_X1 reg_file_reg_30__6_ ( .D(n2588), .CK(clk_i), .Q(reg_file[38]), .QN(
        n3887) );
  DFF_X1 reg_file_reg_29__6_ ( .D(n2589), .CK(clk_i), .Q(reg_file[70]), .QN(
        n3886) );
  DFF_X1 reg_file_reg_28__6_ ( .D(n2590), .CK(clk_i), .Q(reg_file[102]), .QN(
        n4406) );
  DFF_X1 reg_file_reg_27__6_ ( .D(n2591), .CK(clk_i), .Q(reg_file[134]), .QN(
        n4191) );
  DFF_X1 reg_file_reg_2__6_ ( .D(n2616), .CK(clk_i), .Q(reg_file[934]), .QN(
        n4184) );
  DFF_X1 reg_file_reg_1__6_ ( .D(n2617), .CK(clk_i), .Q(reg_file[966]), .QN(
        n4396) );
  DFF_X1 reg_file_reg_0__6_ ( .D(n2618), .CK(clk_i), .Q(reg_file[998]), .QN(
        n3876) );
  DFF_X1 reg_file_reg_31__2_ ( .D(n2715), .CK(clk_i), .Q(reg_file[2]) );
  DFF_X1 reg_file_reg_30__2_ ( .D(n2716), .CK(clk_i), .Q(reg_file[34]) );
  DFF_X1 reg_file_reg_29__2_ ( .D(n2717), .CK(clk_i), .Q(reg_file[66]) );
  DFF_X1 reg_file_reg_28__2_ ( .D(n2718), .CK(clk_i), .Q(reg_file[98]) );
  DFF_X1 reg_file_reg_27__2_ ( .D(n2719), .CK(clk_i), .Q(reg_file[130]) );
  DFF_X1 reg_file_reg_26__2_ ( .D(n2720), .CK(clk_i), .Q(reg_file[162]) );
  DFF_X1 reg_file_reg_25__2_ ( .D(n2721), .CK(clk_i), .Q(reg_file[194]) );
  DFF_X1 reg_file_reg_24__2_ ( .D(n2722), .CK(clk_i), .Q(reg_file[226]) );
  DFF_X1 reg_file_reg_23__2_ ( .D(n2723), .CK(clk_i), .Q(reg_file[258]) );
  DFF_X1 reg_file_reg_22__2_ ( .D(n2724), .CK(clk_i), .Q(reg_file[290]) );
  DFF_X1 reg_file_reg_21__2_ ( .D(n2725), .CK(clk_i), .Q(reg_file[322]) );
  DFF_X1 reg_file_reg_20__2_ ( .D(n2726), .CK(clk_i), .Q(reg_file[354]) );
  DFF_X1 reg_file_reg_19__2_ ( .D(n2727), .CK(clk_i), .Q(reg_file[386]) );
  DFF_X1 reg_file_reg_18__2_ ( .D(n2728), .CK(clk_i), .Q(reg_file[418]) );
  DFF_X1 reg_file_reg_17__2_ ( .D(n2729), .CK(clk_i), .Q(reg_file[450]) );
  DFF_X1 reg_file_reg_16__2_ ( .D(n2730), .CK(clk_i), .Q(reg_file[482]) );
  DFF_X1 reg_file_reg_15__2_ ( .D(n2731), .CK(clk_i), .Q(reg_file[514]) );
  DFF_X1 reg_file_reg_14__2_ ( .D(n2732), .CK(clk_i), .Q(reg_file[546]) );
  DFF_X1 reg_file_reg_13__2_ ( .D(n2733), .CK(clk_i), .Q(reg_file[578]) );
  DFF_X1 reg_file_reg_12__2_ ( .D(n2734), .CK(clk_i), .Q(reg_file[610]) );
  DFF_X1 reg_file_reg_11__2_ ( .D(n2735), .CK(clk_i), .Q(reg_file[642]) );
  DFF_X1 reg_file_reg_10__2_ ( .D(n2736), .CK(clk_i), .Q(reg_file[674]) );
  DFF_X1 reg_file_reg_9__2_ ( .D(n2737), .CK(clk_i), .Q(reg_file[706]) );
  DFF_X1 reg_file_reg_8__2_ ( .D(n2738), .CK(clk_i), .Q(reg_file[738]) );
  DFF_X1 reg_file_reg_7__2_ ( .D(n2739), .CK(clk_i), .Q(reg_file[770]) );
  DFF_X1 reg_file_reg_6__2_ ( .D(n2740), .CK(clk_i), .Q(reg_file[802]) );
  DFF_X1 reg_file_reg_5__2_ ( .D(n2741), .CK(clk_i), .Q(reg_file[834]) );
  DFF_X1 reg_file_reg_4__2_ ( .D(n2742), .CK(clk_i), .Q(reg_file[866]) );
  DFF_X1 reg_file_reg_3__2_ ( .D(n2743), .CK(clk_i), .Q(reg_file[898]) );
  DFF_X1 reg_file_reg_2__2_ ( .D(n2744), .CK(clk_i), .Q(reg_file[930]) );
  DFF_X1 reg_file_reg_1__2_ ( .D(n2745), .CK(clk_i), .Q(reg_file[962]) );
  DFF_X1 reg_file_reg_0__2_ ( .D(n2746), .CK(clk_i), .Q(reg_file[994]) );
  DFF_X1 reg_file_reg_31__29_ ( .D(n1851), .CK(clk_i), .Q(reg_file[29]), .QN(
        n4683) );
  DFF_X1 reg_file_reg_30__29_ ( .D(n1852), .CK(clk_i), .Q(reg_file[61]), .QN(
        n4163) );
  DFF_X1 reg_file_reg_29__29_ ( .D(n1853), .CK(clk_i), .Q(reg_file[93]), .QN(
        n4162) );
  DFF_X1 reg_file_reg_28__29_ ( .D(n1854), .CK(clk_i), .Q(reg_file[125]), .QN(
        n4682) );
  DFF_X1 reg_file_reg_27__29_ ( .D(n1855), .CK(clk_i), .Q(reg_file[157]), .QN(
        n4375) );
  DFF_X1 reg_file_reg_26__29_ ( .D(n1856), .CK(clk_i), .Q(reg_file[189]), .QN(
        n4374) );
  DFF_X1 reg_file_reg_25__29_ ( .D(n1857), .CK(clk_i), .Q(reg_file[221]), .QN(
        n4681) );
  DFF_X1 reg_file_reg_24__29_ ( .D(n1858), .CK(clk_i), .Q(reg_file[253]), .QN(
        n4161) );
  DFF_X1 reg_file_reg_23__29_ ( .D(n1859), .CK(clk_i), .Q(reg_file[285]), .QN(
        n4680) );
  DFF_X1 reg_file_reg_22__29_ ( .D(n1860), .CK(clk_i), .Q(reg_file[317]), .QN(
        n4160) );
  DFF_X1 reg_file_reg_21__29_ ( .D(n1861), .CK(clk_i), .Q(reg_file[349]), .QN(
        n4159) );
  DFF_X1 reg_file_reg_20__29_ ( .D(n1862), .CK(clk_i), .Q(reg_file[381]), .QN(
        n4679) );
  DFF_X1 reg_file_reg_19__29_ ( .D(n1863), .CK(clk_i), .Q(reg_file[413]), .QN(
        n4373) );
  DFF_X1 reg_file_reg_18__29_ ( .D(n1864), .CK(clk_i), .Q(reg_file[445]), .QN(
        n4372) );
  DFF_X1 reg_file_reg_17__29_ ( .D(n1865), .CK(clk_i), .Q(reg_file[477]), .QN(
        n4678) );
  DFF_X1 reg_file_reg_16__29_ ( .D(n1866), .CK(clk_i), .Q(reg_file[509]), .QN(
        n4158) );
  DFF_X1 reg_file_reg_15__29_ ( .D(n1867), .CK(clk_i), .Q(reg_file[541]), .QN(
        n4677) );
  DFF_X1 reg_file_reg_14__29_ ( .D(n1868), .CK(clk_i), .Q(reg_file[573]), .QN(
        n4157) );
  DFF_X1 reg_file_reg_13__29_ ( .D(n1869), .CK(clk_i), .Q(reg_file[605]), .QN(
        n4156) );
  DFF_X1 reg_file_reg_12__29_ ( .D(n1870), .CK(clk_i), .Q(reg_file[637]), .QN(
        n4676) );
  DFF_X1 reg_file_reg_11__29_ ( .D(n1871), .CK(clk_i), .Q(reg_file[669]), .QN(
        n4371) );
  DFF_X1 reg_file_reg_10__29_ ( .D(n1872), .CK(clk_i), .Q(reg_file[701]), .QN(
        n4370) );
  DFF_X1 reg_file_reg_9__29_ ( .D(n1873), .CK(clk_i), .Q(reg_file[733]), .QN(
        n4675) );
  DFF_X1 reg_file_reg_8__29_ ( .D(n1874), .CK(clk_i), .Q(reg_file[765]), .QN(
        n4155) );
  DFF_X1 reg_file_reg_7__29_ ( .D(n1875), .CK(clk_i), .Q(reg_file[797]), .QN(
        n4674) );
  DFF_X1 reg_file_reg_6__29_ ( .D(n1876), .CK(clk_i), .Q(reg_file[829]), .QN(
        n4154) );
  DFF_X1 reg_file_reg_5__29_ ( .D(n1877), .CK(clk_i), .Q(reg_file[861]), .QN(
        n4153) );
  DFF_X1 reg_file_reg_4__29_ ( .D(n1878), .CK(clk_i), .Q(reg_file[893]), .QN(
        n4673) );
  DFF_X1 reg_file_reg_3__29_ ( .D(n1879), .CK(clk_i), .Q(reg_file[925]), .QN(
        n4369) );
  DFF_X1 reg_file_reg_2__29_ ( .D(n1880), .CK(clk_i), .Q(reg_file[957]), .QN(
        n4368) );
  DFF_X1 reg_file_reg_1__29_ ( .D(n1881), .CK(clk_i), .Q(reg_file[989]), .QN(
        n4672) );
  DFF_X1 reg_file_reg_0__29_ ( .D(n1882), .CK(clk_i), .Q(reg_file[1021]), .QN(
        n4152) );
  DFF_X1 reg_file_reg_31__25_ ( .D(n1979), .CK(clk_i), .Q(reg_file[25]), .QN(
        n4635) );
  DFF_X1 reg_file_reg_30__25_ ( .D(n1980), .CK(clk_i), .Q(reg_file[57]), .QN(
        n4115) );
  DFF_X1 reg_file_reg_29__25_ ( .D(n1981), .CK(clk_i), .Q(reg_file[89]), .QN(
        n4114) );
  DFF_X1 reg_file_reg_28__25_ ( .D(n1982), .CK(clk_i), .Q(reg_file[121]), .QN(
        n4634) );
  DFF_X1 reg_file_reg_27__25_ ( .D(n1983), .CK(clk_i), .Q(reg_file[153]), .QN(
        n4343) );
  DFF_X1 reg_file_reg_26__25_ ( .D(n1984), .CK(clk_i), .Q(reg_file[185]), .QN(
        n4342) );
  DFF_X1 reg_file_reg_25__25_ ( .D(n1985), .CK(clk_i), .Q(reg_file[217]), .QN(
        n4633) );
  DFF_X1 reg_file_reg_24__25_ ( .D(n1986), .CK(clk_i), .Q(reg_file[249]), .QN(
        n4113) );
  DFF_X1 reg_file_reg_23__25_ ( .D(n1987), .CK(clk_i), .Q(reg_file[281]), .QN(
        n4632) );
  DFF_X1 reg_file_reg_22__25_ ( .D(n1988), .CK(clk_i), .Q(reg_file[313]), .QN(
        n4112) );
  DFF_X1 reg_file_reg_21__25_ ( .D(n1989), .CK(clk_i), .Q(reg_file[345]), .QN(
        n4111) );
  DFF_X1 reg_file_reg_20__25_ ( .D(n1990), .CK(clk_i), .Q(reg_file[377]), .QN(
        n4631) );
  DFF_X1 reg_file_reg_19__25_ ( .D(n1991), .CK(clk_i), .Q(reg_file[409]), .QN(
        n4341) );
  DFF_X1 reg_file_reg_18__25_ ( .D(n1992), .CK(clk_i), .Q(reg_file[441]), .QN(
        n4340) );
  DFF_X1 reg_file_reg_17__25_ ( .D(n1993), .CK(clk_i), .Q(reg_file[473]), .QN(
        n4630) );
  DFF_X1 reg_file_reg_16__25_ ( .D(n1994), .CK(clk_i), .Q(reg_file[505]), .QN(
        n4110) );
  DFF_X1 reg_file_reg_15__25_ ( .D(n1995), .CK(clk_i), .Q(reg_file[537]), .QN(
        n4629) );
  DFF_X1 reg_file_reg_14__25_ ( .D(n1996), .CK(clk_i), .Q(reg_file[569]), .QN(
        n4109) );
  DFF_X1 reg_file_reg_13__25_ ( .D(n1997), .CK(clk_i), .Q(reg_file[601]), .QN(
        n4108) );
  DFF_X1 reg_file_reg_12__25_ ( .D(n1998), .CK(clk_i), .Q(reg_file[633]), .QN(
        n4628) );
  DFF_X1 reg_file_reg_11__25_ ( .D(n1999), .CK(clk_i), .Q(reg_file[665]), .QN(
        n4339) );
  DFF_X1 reg_file_reg_10__25_ ( .D(n2000), .CK(clk_i), .Q(reg_file[697]), .QN(
        n4338) );
  DFF_X1 reg_file_reg_9__25_ ( .D(n2001), .CK(clk_i), .Q(reg_file[729]), .QN(
        n4627) );
  DFF_X1 reg_file_reg_8__25_ ( .D(n2002), .CK(clk_i), .Q(reg_file[761]), .QN(
        n4107) );
  DFF_X1 reg_file_reg_7__25_ ( .D(n2003), .CK(clk_i), .Q(reg_file[793]), .QN(
        n4626) );
  DFF_X1 reg_file_reg_6__25_ ( .D(n2004), .CK(clk_i), .Q(reg_file[825]), .QN(
        n4106) );
  DFF_X1 reg_file_reg_5__25_ ( .D(n2005), .CK(clk_i), .Q(reg_file[857]), .QN(
        n4105) );
  DFF_X1 reg_file_reg_4__25_ ( .D(n2006), .CK(clk_i), .Q(reg_file[889]), .QN(
        n4625) );
  DFF_X1 reg_file_reg_3__25_ ( .D(n2007), .CK(clk_i), .Q(reg_file[921]), .QN(
        n4337) );
  DFF_X1 reg_file_reg_2__25_ ( .D(n2008), .CK(clk_i), .Q(reg_file[953]), .QN(
        n4336) );
  DFF_X1 reg_file_reg_1__25_ ( .D(n2009), .CK(clk_i), .Q(reg_file[985]), .QN(
        n4624) );
  DFF_X1 reg_file_reg_0__25_ ( .D(n2010), .CK(clk_i), .Q(reg_file[1017]), .QN(
        n4104) );
  DFF_X1 reg_file_reg_31__21_ ( .D(n2107), .CK(clk_i), .Q(reg_file[21]), .QN(
        n4587) );
  DFF_X1 reg_file_reg_30__21_ ( .D(n2108), .CK(clk_i), .Q(reg_file[53]), .QN(
        n4067) );
  DFF_X1 reg_file_reg_29__21_ ( .D(n2109), .CK(clk_i), .Q(reg_file[85]), .QN(
        n4066) );
  DFF_X1 reg_file_reg_28__21_ ( .D(n2110), .CK(clk_i), .Q(reg_file[117]), .QN(
        n4586) );
  DFF_X1 reg_file_reg_27__21_ ( .D(n2111), .CK(clk_i), .Q(reg_file[149]), .QN(
        n4311) );
  DFF_X1 reg_file_reg_26__21_ ( .D(n2112), .CK(clk_i), .Q(reg_file[181]), .QN(
        n4310) );
  DFF_X1 reg_file_reg_25__21_ ( .D(n2113), .CK(clk_i), .Q(reg_file[213]), .QN(
        n4585) );
  DFF_X1 reg_file_reg_24__21_ ( .D(n2114), .CK(clk_i), .Q(reg_file[245]), .QN(
        n4065) );
  DFF_X1 reg_file_reg_23__21_ ( .D(n2115), .CK(clk_i), .Q(reg_file[277]), .QN(
        n4584) );
  DFF_X1 reg_file_reg_22__21_ ( .D(n2116), .CK(clk_i), .Q(reg_file[309]), .QN(
        n4064) );
  DFF_X1 reg_file_reg_21__21_ ( .D(n2117), .CK(clk_i), .Q(reg_file[341]), .QN(
        n4063) );
  DFF_X1 reg_file_reg_20__21_ ( .D(n2118), .CK(clk_i), .Q(reg_file[373]), .QN(
        n4583) );
  DFF_X1 reg_file_reg_19__21_ ( .D(n2119), .CK(clk_i), .Q(reg_file[405]), .QN(
        n4309) );
  DFF_X1 reg_file_reg_18__21_ ( .D(n2120), .CK(clk_i), .Q(reg_file[437]), .QN(
        n4308) );
  DFF_X1 reg_file_reg_17__21_ ( .D(n2121), .CK(clk_i), .Q(reg_file[469]), .QN(
        n4582) );
  DFF_X1 reg_file_reg_16__21_ ( .D(n2122), .CK(clk_i), .Q(reg_file[501]), .QN(
        n4062) );
  DFF_X1 reg_file_reg_15__21_ ( .D(n2123), .CK(clk_i), .Q(reg_file[533]), .QN(
        n4581) );
  DFF_X1 reg_file_reg_14__21_ ( .D(n2124), .CK(clk_i), .Q(reg_file[565]), .QN(
        n4061) );
  DFF_X1 reg_file_reg_13__21_ ( .D(n2125), .CK(clk_i), .Q(reg_file[597]), .QN(
        n4060) );
  DFF_X1 reg_file_reg_12__21_ ( .D(n2126), .CK(clk_i), .Q(reg_file[629]), .QN(
        n4580) );
  DFF_X1 reg_file_reg_11__21_ ( .D(n2127), .CK(clk_i), .Q(reg_file[661]), .QN(
        n4307) );
  DFF_X1 reg_file_reg_10__21_ ( .D(n2128), .CK(clk_i), .Q(reg_file[693]), .QN(
        n4306) );
  DFF_X1 reg_file_reg_9__21_ ( .D(n2129), .CK(clk_i), .Q(reg_file[725]), .QN(
        n4579) );
  DFF_X1 reg_file_reg_8__21_ ( .D(n2130), .CK(clk_i), .Q(reg_file[757]), .QN(
        n4059) );
  DFF_X1 reg_file_reg_7__21_ ( .D(n2131), .CK(clk_i), .Q(reg_file[789]), .QN(
        n4578) );
  DFF_X1 reg_file_reg_6__21_ ( .D(n2132), .CK(clk_i), .Q(reg_file[821]), .QN(
        n4058) );
  DFF_X1 reg_file_reg_5__21_ ( .D(n2133), .CK(clk_i), .Q(reg_file[853]), .QN(
        n4057) );
  DFF_X1 reg_file_reg_4__21_ ( .D(n2134), .CK(clk_i), .Q(reg_file[885]), .QN(
        n4577) );
  DFF_X1 reg_file_reg_3__21_ ( .D(n2135), .CK(clk_i), .Q(reg_file[917]), .QN(
        n4305) );
  DFF_X1 reg_file_reg_2__21_ ( .D(n2136), .CK(clk_i), .Q(reg_file[949]), .QN(
        n4304) );
  DFF_X1 reg_file_reg_1__21_ ( .D(n2137), .CK(clk_i), .Q(reg_file[981]), .QN(
        n4576) );
  DFF_X1 reg_file_reg_0__21_ ( .D(n2138), .CK(clk_i), .Q(reg_file[1013]), .QN(
        n4056) );
  DFF_X1 reg_file_reg_31__17_ ( .D(n2235), .CK(clk_i), .Q(reg_file[17]), .QN(
        n4539) );
  DFF_X1 reg_file_reg_30__17_ ( .D(n2236), .CK(clk_i), .Q(reg_file[49]), .QN(
        n4019) );
  DFF_X1 reg_file_reg_29__17_ ( .D(n2237), .CK(clk_i), .Q(reg_file[81]), .QN(
        n4018) );
  DFF_X1 reg_file_reg_28__17_ ( .D(n2238), .CK(clk_i), .Q(reg_file[113]), .QN(
        n4538) );
  DFF_X1 reg_file_reg_27__17_ ( .D(n2239), .CK(clk_i), .Q(reg_file[145]), .QN(
        n4279) );
  DFF_X1 reg_file_reg_26__17_ ( .D(n2240), .CK(clk_i), .Q(reg_file[177]), .QN(
        n4278) );
  DFF_X1 reg_file_reg_25__17_ ( .D(n2241), .CK(clk_i), .Q(reg_file[209]), .QN(
        n4537) );
  DFF_X1 reg_file_reg_24__17_ ( .D(n2242), .CK(clk_i), .Q(reg_file[241]), .QN(
        n4017) );
  DFF_X1 reg_file_reg_23__17_ ( .D(n2243), .CK(clk_i), .Q(reg_file[273]), .QN(
        n4536) );
  DFF_X1 reg_file_reg_22__17_ ( .D(n2244), .CK(clk_i), .Q(reg_file[305]), .QN(
        n4016) );
  DFF_X1 reg_file_reg_21__17_ ( .D(n2245), .CK(clk_i), .Q(reg_file[337]), .QN(
        n4015) );
  DFF_X1 reg_file_reg_20__17_ ( .D(n2246), .CK(clk_i), .Q(reg_file[369]), .QN(
        n4535) );
  DFF_X1 reg_file_reg_19__17_ ( .D(n2247), .CK(clk_i), .Q(reg_file[401]), .QN(
        n4277) );
  DFF_X1 reg_file_reg_18__17_ ( .D(n2248), .CK(clk_i), .Q(reg_file[433]), .QN(
        n4276) );
  DFF_X1 reg_file_reg_17__17_ ( .D(n2249), .CK(clk_i), .Q(reg_file[465]), .QN(
        n4534) );
  DFF_X1 reg_file_reg_16__17_ ( .D(n2250), .CK(clk_i), .Q(reg_file[497]), .QN(
        n4014) );
  DFF_X1 reg_file_reg_15__17_ ( .D(n2251), .CK(clk_i), .Q(reg_file[529]), .QN(
        n4533) );
  DFF_X1 reg_file_reg_14__17_ ( .D(n2252), .CK(clk_i), .Q(reg_file[561]), .QN(
        n4013) );
  DFF_X1 reg_file_reg_13__17_ ( .D(n2253), .CK(clk_i), .Q(reg_file[593]), .QN(
        n4012) );
  DFF_X1 reg_file_reg_12__17_ ( .D(n2254), .CK(clk_i), .Q(reg_file[625]), .QN(
        n4532) );
  DFF_X1 reg_file_reg_11__17_ ( .D(n2255), .CK(clk_i), .Q(reg_file[657]), .QN(
        n4275) );
  DFF_X1 reg_file_reg_10__17_ ( .D(n2256), .CK(clk_i), .Q(reg_file[689]), .QN(
        n4274) );
  DFF_X1 reg_file_reg_9__17_ ( .D(n2257), .CK(clk_i), .Q(reg_file[721]), .QN(
        n4531) );
  DFF_X1 reg_file_reg_8__17_ ( .D(n2258), .CK(clk_i), .Q(reg_file[753]), .QN(
        n4011) );
  DFF_X1 reg_file_reg_7__17_ ( .D(n2259), .CK(clk_i), .Q(reg_file[785]), .QN(
        n4530) );
  DFF_X1 reg_file_reg_6__17_ ( .D(n2260), .CK(clk_i), .Q(reg_file[817]), .QN(
        n4010) );
  DFF_X1 reg_file_reg_5__17_ ( .D(n2261), .CK(clk_i), .Q(reg_file[849]), .QN(
        n4009) );
  DFF_X1 reg_file_reg_4__17_ ( .D(n2262), .CK(clk_i), .Q(reg_file[881]), .QN(
        n4529) );
  DFF_X1 reg_file_reg_3__17_ ( .D(n2263), .CK(clk_i), .Q(reg_file[913]), .QN(
        n4273) );
  DFF_X1 reg_file_reg_2__17_ ( .D(n2264), .CK(clk_i), .Q(reg_file[945]), .QN(
        n4272) );
  DFF_X1 reg_file_reg_1__17_ ( .D(n2265), .CK(clk_i), .Q(reg_file[977]), .QN(
        n4528) );
  DFF_X1 reg_file_reg_0__17_ ( .D(n2266), .CK(clk_i), .Q(reg_file[1009]), .QN(
        n4008) );
  DFF_X1 reg_file_reg_31__15_ ( .D(n2299), .CK(clk_i), .Q(reg_file[15]), .QN(
        n4515) );
  DFF_X1 reg_file_reg_30__15_ ( .D(n2300), .CK(clk_i), .Q(reg_file[47]), .QN(
        n3995) );
  DFF_X1 reg_file_reg_29__15_ ( .D(n2301), .CK(clk_i), .Q(reg_file[79]), .QN(
        n3994) );
  DFF_X1 reg_file_reg_28__15_ ( .D(n2302), .CK(clk_i), .Q(reg_file[111]), .QN(
        n4514) );
  DFF_X1 reg_file_reg_27__15_ ( .D(n2303), .CK(clk_i), .Q(reg_file[143]), .QN(
        n4263) );
  DFF_X1 reg_file_reg_26__15_ ( .D(n2304), .CK(clk_i), .Q(reg_file[175]), .QN(
        n4262) );
  DFF_X1 reg_file_reg_25__15_ ( .D(n2305), .CK(clk_i), .Q(reg_file[207]), .QN(
        n4513) );
  DFF_X1 reg_file_reg_24__15_ ( .D(n2306), .CK(clk_i), .Q(reg_file[239]), .QN(
        n3993) );
  DFF_X1 reg_file_reg_23__15_ ( .D(n2307), .CK(clk_i), .Q(reg_file[271]), .QN(
        n4512) );
  DFF_X1 reg_file_reg_22__15_ ( .D(n2308), .CK(clk_i), .Q(reg_file[303]), .QN(
        n3992) );
  DFF_X1 reg_file_reg_21__15_ ( .D(n2309), .CK(clk_i), .Q(reg_file[335]), .QN(
        n3991) );
  DFF_X1 reg_file_reg_20__15_ ( .D(n2310), .CK(clk_i), .Q(reg_file[367]), .QN(
        n4511) );
  DFF_X1 reg_file_reg_19__15_ ( .D(n2311), .CK(clk_i), .Q(reg_file[399]), .QN(
        n4261) );
  DFF_X1 reg_file_reg_18__15_ ( .D(n2312), .CK(clk_i), .Q(reg_file[431]), .QN(
        n4260) );
  DFF_X1 reg_file_reg_17__15_ ( .D(n2313), .CK(clk_i), .Q(reg_file[463]), .QN(
        n4510) );
  DFF_X1 reg_file_reg_16__15_ ( .D(n2314), .CK(clk_i), .Q(reg_file[495]), .QN(
        n3990) );
  DFF_X1 reg_file_reg_15__15_ ( .D(n2315), .CK(clk_i), .Q(reg_file[527]), .QN(
        n4509) );
  DFF_X1 reg_file_reg_14__15_ ( .D(n2316), .CK(clk_i), .Q(reg_file[559]), .QN(
        n3989) );
  DFF_X1 reg_file_reg_13__15_ ( .D(n2317), .CK(clk_i), .Q(reg_file[591]), .QN(
        n3988) );
  DFF_X1 reg_file_reg_12__15_ ( .D(n2318), .CK(clk_i), .Q(reg_file[623]), .QN(
        n4508) );
  DFF_X1 reg_file_reg_11__15_ ( .D(n2319), .CK(clk_i), .Q(reg_file[655]), .QN(
        n4259) );
  DFF_X1 reg_file_reg_10__15_ ( .D(n2320), .CK(clk_i), .Q(reg_file[687]), .QN(
        n4258) );
  DFF_X1 reg_file_reg_9__15_ ( .D(n2321), .CK(clk_i), .Q(reg_file[719]), .QN(
        n4507) );
  DFF_X1 reg_file_reg_8__15_ ( .D(n2322), .CK(clk_i), .Q(reg_file[751]), .QN(
        n3987) );
  DFF_X1 reg_file_reg_7__15_ ( .D(n2323), .CK(clk_i), .Q(reg_file[783]), .QN(
        n4506) );
  DFF_X1 reg_file_reg_6__15_ ( .D(n2324), .CK(clk_i), .Q(reg_file[815]), .QN(
        n3986) );
  DFF_X1 reg_file_reg_5__15_ ( .D(n2325), .CK(clk_i), .Q(reg_file[847]), .QN(
        n3985) );
  DFF_X1 reg_file_reg_4__15_ ( .D(n2326), .CK(clk_i), .Q(reg_file[879]), .QN(
        n4505) );
  DFF_X1 reg_file_reg_3__15_ ( .D(n2327), .CK(clk_i), .Q(reg_file[911]), .QN(
        n4257) );
  DFF_X1 reg_file_reg_2__15_ ( .D(n2328), .CK(clk_i), .Q(reg_file[943]), .QN(
        n4256) );
  DFF_X1 reg_file_reg_1__15_ ( .D(n2329), .CK(clk_i), .Q(reg_file[975]), .QN(
        n4504) );
  DFF_X1 reg_file_reg_0__15_ ( .D(n2330), .CK(clk_i), .Q(reg_file[1007]), .QN(
        n3984) );
  DFF_X1 reg_file_reg_31__11_ ( .D(n2427), .CK(clk_i), .Q(reg_file[11]), .QN(
        n4467) );
  DFF_X1 reg_file_reg_30__11_ ( .D(n2428), .CK(clk_i), .Q(reg_file[43]), .QN(
        n3947) );
  DFF_X1 reg_file_reg_29__11_ ( .D(n2429), .CK(clk_i), .Q(reg_file[75]), .QN(
        n3946) );
  DFF_X1 reg_file_reg_28__11_ ( .D(n2430), .CK(clk_i), .Q(reg_file[107]), .QN(
        n4466) );
  DFF_X1 reg_file_reg_27__11_ ( .D(n2431), .CK(clk_i), .Q(reg_file[139]), .QN(
        n4231) );
  DFF_X1 reg_file_reg_26__11_ ( .D(n2432), .CK(clk_i), .Q(reg_file[171]), .QN(
        n4230) );
  DFF_X1 reg_file_reg_25__11_ ( .D(n2433), .CK(clk_i), .Q(reg_file[203]), .QN(
        n4465) );
  DFF_X1 reg_file_reg_24__11_ ( .D(n2434), .CK(clk_i), .Q(reg_file[235]), .QN(
        n3945) );
  DFF_X1 reg_file_reg_23__11_ ( .D(n2435), .CK(clk_i), .Q(reg_file[267]), .QN(
        n4464) );
  DFF_X1 reg_file_reg_22__11_ ( .D(n2436), .CK(clk_i), .Q(reg_file[299]), .QN(
        n3944) );
  DFF_X1 reg_file_reg_21__11_ ( .D(n2437), .CK(clk_i), .Q(reg_file[331]), .QN(
        n3943) );
  DFF_X1 reg_file_reg_20__11_ ( .D(n2438), .CK(clk_i), .Q(reg_file[363]), .QN(
        n4463) );
  DFF_X1 reg_file_reg_19__11_ ( .D(n2439), .CK(clk_i), .Q(reg_file[395]), .QN(
        n4229) );
  DFF_X1 reg_file_reg_18__11_ ( .D(n2440), .CK(clk_i), .Q(reg_file[427]), .QN(
        n4228) );
  DFF_X1 reg_file_reg_17__11_ ( .D(n2441), .CK(clk_i), .Q(reg_file[459]), .QN(
        n4462) );
  DFF_X1 reg_file_reg_16__11_ ( .D(n2442), .CK(clk_i), .Q(reg_file[491]), .QN(
        n3942) );
  DFF_X1 reg_file_reg_15__11_ ( .D(n2443), .CK(clk_i), .Q(reg_file[523]), .QN(
        n4461) );
  DFF_X1 reg_file_reg_14__11_ ( .D(n2444), .CK(clk_i), .Q(reg_file[555]), .QN(
        n3941) );
  DFF_X1 reg_file_reg_13__11_ ( .D(n2445), .CK(clk_i), .Q(reg_file[587]), .QN(
        n3940) );
  DFF_X1 reg_file_reg_12__11_ ( .D(n2446), .CK(clk_i), .Q(reg_file[619]), .QN(
        n4460) );
  DFF_X1 reg_file_reg_11__11_ ( .D(n2447), .CK(clk_i), .Q(reg_file[651]), .QN(
        n4227) );
  DFF_X1 reg_file_reg_10__11_ ( .D(n2448), .CK(clk_i), .Q(reg_file[683]), .QN(
        n4226) );
  DFF_X1 reg_file_reg_9__11_ ( .D(n2449), .CK(clk_i), .Q(reg_file[715]), .QN(
        n4459) );
  DFF_X1 reg_file_reg_8__11_ ( .D(n2450), .CK(clk_i), .Q(reg_file[747]), .QN(
        n3939) );
  DFF_X1 reg_file_reg_7__11_ ( .D(n2451), .CK(clk_i), .Q(reg_file[779]), .QN(
        n4458) );
  DFF_X1 reg_file_reg_6__11_ ( .D(n2452), .CK(clk_i), .Q(reg_file[811]), .QN(
        n3938) );
  DFF_X1 reg_file_reg_5__11_ ( .D(n2453), .CK(clk_i), .Q(reg_file[843]), .QN(
        n3937) );
  DFF_X1 reg_file_reg_4__11_ ( .D(n2454), .CK(clk_i), .Q(reg_file[875]), .QN(
        n4457) );
  DFF_X1 reg_file_reg_3__11_ ( .D(n2455), .CK(clk_i), .Q(reg_file[907]), .QN(
        n4225) );
  DFF_X1 reg_file_reg_2__11_ ( .D(n2456), .CK(clk_i), .Q(reg_file[939]), .QN(
        n4224) );
  DFF_X1 reg_file_reg_1__11_ ( .D(n2457), .CK(clk_i), .Q(reg_file[971]), .QN(
        n4456) );
  DFF_X1 reg_file_reg_0__11_ ( .D(n2458), .CK(clk_i), .Q(reg_file[1003]), .QN(
        n3936) );
  DFF_X1 reg_file_reg_31__3_ ( .D(n2683), .CK(clk_i), .Q(reg_file[3]) );
  DFF_X1 reg_file_reg_30__3_ ( .D(n2684), .CK(clk_i), .Q(reg_file[35]) );
  DFF_X1 reg_file_reg_29__3_ ( .D(n2685), .CK(clk_i), .Q(reg_file[67]) );
  DFF_X1 reg_file_reg_28__3_ ( .D(n2686), .CK(clk_i), .Q(reg_file[99]) );
  DFF_X1 reg_file_reg_27__3_ ( .D(n2687), .CK(clk_i), .Q(reg_file[131]) );
  DFF_X1 reg_file_reg_26__3_ ( .D(n2688), .CK(clk_i), .Q(reg_file[163]) );
  DFF_X1 reg_file_reg_25__3_ ( .D(n2689), .CK(clk_i), .Q(reg_file[195]) );
  DFF_X1 reg_file_reg_24__3_ ( .D(n2690), .CK(clk_i), .Q(reg_file[227]) );
  DFF_X1 reg_file_reg_23__3_ ( .D(n2691), .CK(clk_i), .Q(reg_file[259]) );
  DFF_X1 reg_file_reg_22__3_ ( .D(n2692), .CK(clk_i), .Q(reg_file[291]) );
  DFF_X1 reg_file_reg_21__3_ ( .D(n2693), .CK(clk_i), .Q(reg_file[323]) );
  DFF_X1 reg_file_reg_20__3_ ( .D(n2694), .CK(clk_i), .Q(reg_file[355]) );
  DFF_X1 reg_file_reg_19__3_ ( .D(n2695), .CK(clk_i), .Q(reg_file[387]) );
  DFF_X1 reg_file_reg_18__3_ ( .D(n2696), .CK(clk_i), .Q(reg_file[419]) );
  DFF_X1 reg_file_reg_17__3_ ( .D(n2697), .CK(clk_i), .Q(reg_file[451]) );
  DFF_X1 reg_file_reg_16__3_ ( .D(n2698), .CK(clk_i), .Q(reg_file[483]) );
  DFF_X1 reg_file_reg_15__3_ ( .D(n2699), .CK(clk_i), .Q(reg_file[515]) );
  DFF_X1 reg_file_reg_14__3_ ( .D(n2700), .CK(clk_i), .Q(reg_file[547]) );
  DFF_X1 reg_file_reg_13__3_ ( .D(n2701), .CK(clk_i), .Q(reg_file[579]) );
  DFF_X1 reg_file_reg_12__3_ ( .D(n2702), .CK(clk_i), .Q(reg_file[611]) );
  DFF_X1 reg_file_reg_11__3_ ( .D(n2703), .CK(clk_i), .Q(reg_file[643]) );
  DFF_X1 reg_file_reg_10__3_ ( .D(n2704), .CK(clk_i), .Q(reg_file[675]) );
  DFF_X1 reg_file_reg_9__3_ ( .D(n2705), .CK(clk_i), .Q(reg_file[707]) );
  DFF_X1 reg_file_reg_8__3_ ( .D(n2706), .CK(clk_i), .Q(reg_file[739]) );
  DFF_X1 reg_file_reg_7__3_ ( .D(n2707), .CK(clk_i), .Q(reg_file[771]) );
  DFF_X1 reg_file_reg_6__3_ ( .D(n2708), .CK(clk_i), .Q(reg_file[803]) );
  DFF_X1 reg_file_reg_5__3_ ( .D(n2709), .CK(clk_i), .Q(reg_file[835]) );
  DFF_X1 reg_file_reg_4__3_ ( .D(n2710), .CK(clk_i), .Q(reg_file[867]) );
  DFF_X1 reg_file_reg_3__3_ ( .D(n2711), .CK(clk_i), .Q(reg_file[899]) );
  DFF_X1 reg_file_reg_2__3_ ( .D(n2712), .CK(clk_i), .Q(reg_file[931]) );
  DFF_X1 reg_file_reg_1__3_ ( .D(n2713), .CK(clk_i), .Q(reg_file[963]) );
  DFF_X1 reg_file_reg_0__3_ ( .D(n2714), .CK(clk_i), .Q(reg_file[995]) );
  DFF_X1 reg_file_reg_31__28_ ( .D(n1883), .CK(clk_i), .Q(reg_file[28]), .QN(
        n4671) );
  DFF_X1 reg_file_reg_30__28_ ( .D(n1884), .CK(clk_i), .Q(reg_file[60]), .QN(
        n4151) );
  DFF_X1 reg_file_reg_29__28_ ( .D(n1885), .CK(clk_i), .Q(reg_file[92]), .QN(
        n4150) );
  DFF_X1 reg_file_reg_28__28_ ( .D(n1886), .CK(clk_i), .Q(reg_file[124]), .QN(
        n4670) );
  DFF_X1 reg_file_reg_27__28_ ( .D(n1887), .CK(clk_i), .Q(reg_file[156]), .QN(
        n4367) );
  DFF_X1 reg_file_reg_26__28_ ( .D(n1888), .CK(clk_i), .Q(reg_file[188]), .QN(
        n4366) );
  DFF_X1 reg_file_reg_25__28_ ( .D(n1889), .CK(clk_i), .Q(reg_file[220]), .QN(
        n4669) );
  DFF_X1 reg_file_reg_24__28_ ( .D(n1890), .CK(clk_i), .Q(reg_file[252]), .QN(
        n4149) );
  DFF_X1 reg_file_reg_23__28_ ( .D(n1891), .CK(clk_i), .Q(reg_file[284]), .QN(
        n4668) );
  DFF_X1 reg_file_reg_22__28_ ( .D(n1892), .CK(clk_i), .Q(reg_file[316]), .QN(
        n4148) );
  DFF_X1 reg_file_reg_21__28_ ( .D(n1893), .CK(clk_i), .Q(reg_file[348]), .QN(
        n4147) );
  DFF_X1 reg_file_reg_20__28_ ( .D(n1894), .CK(clk_i), .Q(reg_file[380]), .QN(
        n4667) );
  DFF_X1 reg_file_reg_19__28_ ( .D(n1895), .CK(clk_i), .Q(reg_file[412]), .QN(
        n4365) );
  DFF_X1 reg_file_reg_18__28_ ( .D(n1896), .CK(clk_i), .Q(reg_file[444]), .QN(
        n4364) );
  DFF_X1 reg_file_reg_17__28_ ( .D(n1897), .CK(clk_i), .Q(reg_file[476]), .QN(
        n4666) );
  DFF_X1 reg_file_reg_16__28_ ( .D(n1898), .CK(clk_i), .Q(reg_file[508]), .QN(
        n4146) );
  DFF_X1 reg_file_reg_15__28_ ( .D(n1899), .CK(clk_i), .Q(reg_file[540]), .QN(
        n4665) );
  DFF_X1 reg_file_reg_14__28_ ( .D(n1900), .CK(clk_i), .Q(reg_file[572]), .QN(
        n4145) );
  DFF_X1 reg_file_reg_13__28_ ( .D(n1901), .CK(clk_i), .Q(reg_file[604]), .QN(
        n4144) );
  DFF_X1 reg_file_reg_12__28_ ( .D(n1902), .CK(clk_i), .Q(reg_file[636]), .QN(
        n4664) );
  DFF_X1 reg_file_reg_11__28_ ( .D(n1903), .CK(clk_i), .Q(reg_file[668]), .QN(
        n4363) );
  DFF_X1 reg_file_reg_10__28_ ( .D(n1904), .CK(clk_i), .Q(reg_file[700]), .QN(
        n4362) );
  DFF_X1 reg_file_reg_9__28_ ( .D(n1905), .CK(clk_i), .Q(reg_file[732]), .QN(
        n4663) );
  DFF_X1 reg_file_reg_8__28_ ( .D(n1906), .CK(clk_i), .Q(reg_file[764]), .QN(
        n4143) );
  DFF_X1 reg_file_reg_7__28_ ( .D(n1907), .CK(clk_i), .Q(reg_file[796]), .QN(
        n4662) );
  DFF_X1 reg_file_reg_6__28_ ( .D(n1908), .CK(clk_i), .Q(reg_file[828]), .QN(
        n4142) );
  DFF_X1 reg_file_reg_5__28_ ( .D(n1909), .CK(clk_i), .Q(reg_file[860]), .QN(
        n4141) );
  DFF_X1 reg_file_reg_4__28_ ( .D(n1910), .CK(clk_i), .Q(reg_file[892]), .QN(
        n4661) );
  DFF_X1 reg_file_reg_3__28_ ( .D(n1911), .CK(clk_i), .Q(reg_file[924]), .QN(
        n4361) );
  DFF_X1 reg_file_reg_2__28_ ( .D(n1912), .CK(clk_i), .Q(reg_file[956]), .QN(
        n4360) );
  DFF_X1 reg_file_reg_1__28_ ( .D(n1913), .CK(clk_i), .Q(reg_file[988]), .QN(
        n4660) );
  DFF_X1 reg_file_reg_0__28_ ( .D(n1914), .CK(clk_i), .Q(reg_file[1020]), .QN(
        n4140) );
  DFF_X1 reg_file_reg_31__24_ ( .D(n2011), .CK(clk_i), .Q(reg_file[24]), .QN(
        n4623) );
  DFF_X1 reg_file_reg_30__24_ ( .D(n2012), .CK(clk_i), .Q(reg_file[56]), .QN(
        n4103) );
  DFF_X1 reg_file_reg_29__24_ ( .D(n2013), .CK(clk_i), .Q(reg_file[88]), .QN(
        n4102) );
  DFF_X1 reg_file_reg_28__24_ ( .D(n2014), .CK(clk_i), .Q(reg_file[120]), .QN(
        n4622) );
  DFF_X1 reg_file_reg_27__24_ ( .D(n2015), .CK(clk_i), .Q(reg_file[152]), .QN(
        n4335) );
  DFF_X1 reg_file_reg_26__24_ ( .D(n2016), .CK(clk_i), .Q(reg_file[184]), .QN(
        n4334) );
  DFF_X1 reg_file_reg_25__24_ ( .D(n2017), .CK(clk_i), .Q(reg_file[216]), .QN(
        n4621) );
  DFF_X1 reg_file_reg_24__24_ ( .D(n2018), .CK(clk_i), .Q(reg_file[248]), .QN(
        n4101) );
  DFF_X1 reg_file_reg_23__24_ ( .D(n2019), .CK(clk_i), .Q(reg_file[280]), .QN(
        n4620) );
  DFF_X1 reg_file_reg_22__24_ ( .D(n2020), .CK(clk_i), .Q(reg_file[312]), .QN(
        n4100) );
  DFF_X1 reg_file_reg_21__24_ ( .D(n2021), .CK(clk_i), .Q(reg_file[344]), .QN(
        n4099) );
  DFF_X1 reg_file_reg_20__24_ ( .D(n2022), .CK(clk_i), .Q(reg_file[376]), .QN(
        n4619) );
  DFF_X1 reg_file_reg_19__24_ ( .D(n2023), .CK(clk_i), .Q(reg_file[408]), .QN(
        n4333) );
  DFF_X1 reg_file_reg_18__24_ ( .D(n2024), .CK(clk_i), .Q(reg_file[440]), .QN(
        n4332) );
  DFF_X1 reg_file_reg_17__24_ ( .D(n2025), .CK(clk_i), .Q(reg_file[472]), .QN(
        n4618) );
  DFF_X1 reg_file_reg_16__24_ ( .D(n2026), .CK(clk_i), .Q(reg_file[504]), .QN(
        n4098) );
  DFF_X1 reg_file_reg_15__24_ ( .D(n2027), .CK(clk_i), .Q(reg_file[536]), .QN(
        n4617) );
  DFF_X1 reg_file_reg_14__24_ ( .D(n2028), .CK(clk_i), .Q(reg_file[568]), .QN(
        n4097) );
  DFF_X1 reg_file_reg_13__24_ ( .D(n2029), .CK(clk_i), .Q(reg_file[600]), .QN(
        n4096) );
  DFF_X1 reg_file_reg_12__24_ ( .D(n2030), .CK(clk_i), .Q(reg_file[632]), .QN(
        n4616) );
  DFF_X1 reg_file_reg_11__24_ ( .D(n2031), .CK(clk_i), .Q(reg_file[664]), .QN(
        n4331) );
  DFF_X1 reg_file_reg_10__24_ ( .D(n2032), .CK(clk_i), .Q(reg_file[696]), .QN(
        n4330) );
  DFF_X1 reg_file_reg_9__24_ ( .D(n2033), .CK(clk_i), .Q(reg_file[728]), .QN(
        n4615) );
  DFF_X1 reg_file_reg_8__24_ ( .D(n2034), .CK(clk_i), .Q(reg_file[760]), .QN(
        n4095) );
  DFF_X1 reg_file_reg_7__24_ ( .D(n2035), .CK(clk_i), .Q(reg_file[792]), .QN(
        n4614) );
  DFF_X1 reg_file_reg_6__24_ ( .D(n2036), .CK(clk_i), .Q(reg_file[824]), .QN(
        n4094) );
  DFF_X1 reg_file_reg_5__24_ ( .D(n2037), .CK(clk_i), .Q(reg_file[856]), .QN(
        n4093) );
  DFF_X1 reg_file_reg_4__24_ ( .D(n2038), .CK(clk_i), .Q(reg_file[888]), .QN(
        n4613) );
  DFF_X1 reg_file_reg_3__24_ ( .D(n2039), .CK(clk_i), .Q(reg_file[920]), .QN(
        n4329) );
  DFF_X1 reg_file_reg_2__24_ ( .D(n2040), .CK(clk_i), .Q(reg_file[952]), .QN(
        n4328) );
  DFF_X1 reg_file_reg_1__24_ ( .D(n2041), .CK(clk_i), .Q(reg_file[984]), .QN(
        n4612) );
  DFF_X1 reg_file_reg_0__24_ ( .D(n2042), .CK(clk_i), .Q(reg_file[1016]), .QN(
        n4092) );
  DFF_X1 reg_file_reg_31__20_ ( .D(n2139), .CK(clk_i), .Q(reg_file[20]), .QN(
        n4575) );
  DFF_X1 reg_file_reg_30__20_ ( .D(n2140), .CK(clk_i), .Q(reg_file[52]), .QN(
        n4055) );
  DFF_X1 reg_file_reg_29__20_ ( .D(n2141), .CK(clk_i), .Q(reg_file[84]), .QN(
        n4054) );
  DFF_X1 reg_file_reg_28__20_ ( .D(n2142), .CK(clk_i), .Q(reg_file[116]), .QN(
        n4574) );
  DFF_X1 reg_file_reg_27__20_ ( .D(n2143), .CK(clk_i), .Q(reg_file[148]), .QN(
        n4303) );
  DFF_X1 reg_file_reg_26__20_ ( .D(n2144), .CK(clk_i), .Q(reg_file[180]), .QN(
        n4302) );
  DFF_X1 reg_file_reg_25__20_ ( .D(n2145), .CK(clk_i), .Q(reg_file[212]), .QN(
        n4573) );
  DFF_X1 reg_file_reg_24__20_ ( .D(n2146), .CK(clk_i), .Q(reg_file[244]), .QN(
        n4053) );
  DFF_X1 reg_file_reg_23__20_ ( .D(n2147), .CK(clk_i), .Q(reg_file[276]), .QN(
        n4572) );
  DFF_X1 reg_file_reg_22__20_ ( .D(n2148), .CK(clk_i), .Q(reg_file[308]), .QN(
        n4052) );
  DFF_X1 reg_file_reg_21__20_ ( .D(n2149), .CK(clk_i), .Q(reg_file[340]), .QN(
        n4051) );
  DFF_X1 reg_file_reg_20__20_ ( .D(n2150), .CK(clk_i), .Q(reg_file[372]), .QN(
        n4571) );
  DFF_X1 reg_file_reg_19__20_ ( .D(n2151), .CK(clk_i), .Q(reg_file[404]), .QN(
        n4301) );
  DFF_X1 reg_file_reg_18__20_ ( .D(n2152), .CK(clk_i), .Q(reg_file[436]), .QN(
        n4300) );
  DFF_X1 reg_file_reg_17__20_ ( .D(n2153), .CK(clk_i), .Q(reg_file[468]), .QN(
        n4570) );
  DFF_X1 reg_file_reg_16__20_ ( .D(n2154), .CK(clk_i), .Q(reg_file[500]), .QN(
        n4050) );
  DFF_X1 reg_file_reg_15__20_ ( .D(n2155), .CK(clk_i), .Q(reg_file[532]), .QN(
        n4569) );
  DFF_X1 reg_file_reg_14__20_ ( .D(n2156), .CK(clk_i), .Q(reg_file[564]), .QN(
        n4049) );
  DFF_X1 reg_file_reg_13__20_ ( .D(n2157), .CK(clk_i), .Q(reg_file[596]), .QN(
        n4048) );
  DFF_X1 reg_file_reg_12__20_ ( .D(n2158), .CK(clk_i), .Q(reg_file[628]), .QN(
        n4568) );
  DFF_X1 reg_file_reg_11__20_ ( .D(n2159), .CK(clk_i), .Q(reg_file[660]), .QN(
        n4299) );
  DFF_X1 reg_file_reg_10__20_ ( .D(n2160), .CK(clk_i), .Q(reg_file[692]), .QN(
        n4298) );
  DFF_X1 reg_file_reg_9__20_ ( .D(n2161), .CK(clk_i), .Q(reg_file[724]), .QN(
        n4567) );
  DFF_X1 reg_file_reg_8__20_ ( .D(n2162), .CK(clk_i), .Q(reg_file[756]), .QN(
        n4047) );
  DFF_X1 reg_file_reg_7__20_ ( .D(n2163), .CK(clk_i), .Q(reg_file[788]), .QN(
        n4566) );
  DFF_X1 reg_file_reg_6__20_ ( .D(n2164), .CK(clk_i), .Q(reg_file[820]), .QN(
        n4046) );
  DFF_X1 reg_file_reg_5__20_ ( .D(n2165), .CK(clk_i), .Q(reg_file[852]), .QN(
        n4045) );
  DFF_X1 reg_file_reg_4__20_ ( .D(n2166), .CK(clk_i), .Q(reg_file[884]), .QN(
        n4565) );
  DFF_X1 reg_file_reg_3__20_ ( .D(n2167), .CK(clk_i), .Q(reg_file[916]), .QN(
        n4297) );
  DFF_X1 reg_file_reg_2__20_ ( .D(n2168), .CK(clk_i), .Q(reg_file[948]), .QN(
        n4296) );
  DFF_X1 reg_file_reg_1__20_ ( .D(n2169), .CK(clk_i), .Q(reg_file[980]), .QN(
        n4564) );
  DFF_X1 reg_file_reg_0__20_ ( .D(n2170), .CK(clk_i), .Q(reg_file[1012]), .QN(
        n4044) );
  DFF_X1 reg_file_reg_31__0_ ( .D(n1755), .CK(clk_i), .Q(reg_file[0]) );
  DFF_X1 reg_file_reg_30__0_ ( .D(n1756), .CK(clk_i), .Q(reg_file[32]) );
  DFF_X1 reg_file_reg_29__0_ ( .D(n1757), .CK(clk_i), .Q(reg_file[64]) );
  DFF_X1 reg_file_reg_28__0_ ( .D(n1758), .CK(clk_i), .Q(reg_file[96]) );
  DFF_X1 reg_file_reg_27__0_ ( .D(n1759), .CK(clk_i), .Q(reg_file[128]) );
  DFF_X1 reg_file_reg_26__0_ ( .D(n1760), .CK(clk_i), .Q(reg_file[160]) );
  DFF_X1 reg_file_reg_25__0_ ( .D(n1761), .CK(clk_i), .Q(reg_file[192]) );
  DFF_X1 reg_file_reg_24__0_ ( .D(n1762), .CK(clk_i), .Q(reg_file[224]) );
  DFF_X1 reg_file_reg_23__0_ ( .D(n1763), .CK(clk_i), .Q(reg_file[256]) );
  DFF_X1 reg_file_reg_22__0_ ( .D(n1764), .CK(clk_i), .Q(reg_file[288]) );
  DFF_X1 reg_file_reg_21__0_ ( .D(n1765), .CK(clk_i), .Q(reg_file[320]) );
  DFF_X1 reg_file_reg_20__0_ ( .D(n1766), .CK(clk_i), .Q(reg_file[352]) );
  DFF_X1 reg_file_reg_19__0_ ( .D(n1767), .CK(clk_i), .Q(reg_file[384]) );
  DFF_X1 reg_file_reg_18__0_ ( .D(n1768), .CK(clk_i), .Q(reg_file[416]) );
  DFF_X1 reg_file_reg_17__0_ ( .D(n1769), .CK(clk_i), .Q(reg_file[448]) );
  DFF_X1 reg_file_reg_16__0_ ( .D(n1770), .CK(clk_i), .Q(reg_file[480]) );
  DFF_X1 reg_file_reg_15__0_ ( .D(n1771), .CK(clk_i), .Q(reg_file[512]) );
  DFF_X1 reg_file_reg_14__0_ ( .D(n1772), .CK(clk_i), .Q(reg_file[544]) );
  DFF_X1 reg_file_reg_13__0_ ( .D(n1773), .CK(clk_i), .Q(reg_file[576]) );
  DFF_X1 reg_file_reg_12__0_ ( .D(n1774), .CK(clk_i), .Q(reg_file[608]) );
  DFF_X1 reg_file_reg_11__0_ ( .D(n1775), .CK(clk_i), .Q(reg_file[640]) );
  DFF_X1 reg_file_reg_10__0_ ( .D(n1776), .CK(clk_i), .Q(reg_file[672]) );
  DFF_X1 reg_file_reg_9__0_ ( .D(n1777), .CK(clk_i), .Q(reg_file[704]) );
  DFF_X1 reg_file_reg_8__0_ ( .D(n1778), .CK(clk_i), .Q(reg_file[736]) );
  DFF_X1 reg_file_reg_7__0_ ( .D(n1779), .CK(clk_i), .Q(reg_file[768]) );
  DFF_X1 reg_file_reg_6__0_ ( .D(n1780), .CK(clk_i), .Q(reg_file[800]) );
  DFF_X1 reg_file_reg_5__0_ ( .D(n1781), .CK(clk_i), .Q(reg_file[832]) );
  DFF_X1 reg_file_reg_4__0_ ( .D(n1782), .CK(clk_i), .Q(reg_file[864]) );
  DFF_X1 reg_file_reg_3__0_ ( .D(n1783), .CK(clk_i), .Q(reg_file[896]) );
  DFF_X1 reg_file_reg_2__0_ ( .D(n1784), .CK(clk_i), .Q(reg_file[928]) );
  DFF_X1 reg_file_reg_1__0_ ( .D(n1785), .CK(clk_i), .Q(reg_file[960]) );
  DFF_X1 reg_file_reg_0__0_ ( .D(n1786), .CK(clk_i), .Q(reg_file[992]) );
  DFF_X1 reg_file_reg_31__12_ ( .D(n2395), .CK(clk_i), .Q(reg_file[12]), .QN(
        n4479) );
  DFF_X1 reg_file_reg_30__12_ ( .D(n2396), .CK(clk_i), .Q(reg_file[44]), .QN(
        n3959) );
  DFF_X1 reg_file_reg_29__12_ ( .D(n2397), .CK(clk_i), .Q(reg_file[76]), .QN(
        n3958) );
  DFF_X1 reg_file_reg_28__12_ ( .D(n2398), .CK(clk_i), .Q(reg_file[108]), .QN(
        n4478) );
  DFF_X1 reg_file_reg_27__12_ ( .D(n2399), .CK(clk_i), .Q(reg_file[140]), .QN(
        n4239) );
  DFF_X1 reg_file_reg_26__12_ ( .D(n2400), .CK(clk_i), .Q(reg_file[172]), .QN(
        n4238) );
  DFF_X1 reg_file_reg_25__12_ ( .D(n2401), .CK(clk_i), .Q(reg_file[204]), .QN(
        n4477) );
  DFF_X1 reg_file_reg_24__12_ ( .D(n2402), .CK(clk_i), .Q(reg_file[236]), .QN(
        n3957) );
  DFF_X1 reg_file_reg_23__12_ ( .D(n2403), .CK(clk_i), .Q(reg_file[268]), .QN(
        n4476) );
  DFF_X1 reg_file_reg_22__12_ ( .D(n2404), .CK(clk_i), .Q(reg_file[300]), .QN(
        n3956) );
  DFF_X1 reg_file_reg_21__12_ ( .D(n2405), .CK(clk_i), .Q(reg_file[332]), .QN(
        n3955) );
  DFF_X1 reg_file_reg_20__12_ ( .D(n2406), .CK(clk_i), .Q(reg_file[364]), .QN(
        n4475) );
  DFF_X1 reg_file_reg_19__12_ ( .D(n2407), .CK(clk_i), .Q(reg_file[396]), .QN(
        n4237) );
  DFF_X1 reg_file_reg_18__12_ ( .D(n2408), .CK(clk_i), .Q(reg_file[428]), .QN(
        n4236) );
  DFF_X1 reg_file_reg_17__12_ ( .D(n2409), .CK(clk_i), .Q(reg_file[460]), .QN(
        n4474) );
  DFF_X1 reg_file_reg_16__12_ ( .D(n2410), .CK(clk_i), .Q(reg_file[492]), .QN(
        n3954) );
  DFF_X1 reg_file_reg_15__12_ ( .D(n2411), .CK(clk_i), .Q(reg_file[524]), .QN(
        n4473) );
  DFF_X1 reg_file_reg_14__12_ ( .D(n2412), .CK(clk_i), .Q(reg_file[556]), .QN(
        n3953) );
  DFF_X1 reg_file_reg_13__12_ ( .D(n2413), .CK(clk_i), .Q(reg_file[588]), .QN(
        n3952) );
  DFF_X1 reg_file_reg_12__12_ ( .D(n2414), .CK(clk_i), .Q(reg_file[620]), .QN(
        n4472) );
  DFF_X1 reg_file_reg_11__12_ ( .D(n2415), .CK(clk_i), .Q(reg_file[652]), .QN(
        n4235) );
  DFF_X1 reg_file_reg_10__12_ ( .D(n2416), .CK(clk_i), .Q(reg_file[684]), .QN(
        n4234) );
  DFF_X1 reg_file_reg_9__12_ ( .D(n2417), .CK(clk_i), .Q(reg_file[716]), .QN(
        n4471) );
  DFF_X1 reg_file_reg_8__12_ ( .D(n2418), .CK(clk_i), .Q(reg_file[748]), .QN(
        n3951) );
  DFF_X1 reg_file_reg_7__12_ ( .D(n2419), .CK(clk_i), .Q(reg_file[780]), .QN(
        n4470) );
  DFF_X1 reg_file_reg_6__12_ ( .D(n2420), .CK(clk_i), .Q(reg_file[812]), .QN(
        n3950) );
  DFF_X1 reg_file_reg_5__12_ ( .D(n2421), .CK(clk_i), .Q(reg_file[844]), .QN(
        n3949) );
  DFF_X1 reg_file_reg_4__12_ ( .D(n2422), .CK(clk_i), .Q(reg_file[876]), .QN(
        n4469) );
  DFF_X1 reg_file_reg_3__12_ ( .D(n2423), .CK(clk_i), .Q(reg_file[908]), .QN(
        n4233) );
  DFF_X1 reg_file_reg_2__12_ ( .D(n2424), .CK(clk_i), .Q(reg_file[940]), .QN(
        n4232) );
  DFF_X1 reg_file_reg_1__12_ ( .D(n2425), .CK(clk_i), .Q(reg_file[972]), .QN(
        n4468) );
  DFF_X1 reg_file_reg_0__12_ ( .D(n2426), .CK(clk_i), .Q(reg_file[1004]), .QN(
        n3948) );
  DFF_X1 reg_file_reg_31__8_ ( .D(n2523), .CK(clk_i), .Q(reg_file[8]), .QN(
        n4431) );
  DFF_X1 reg_file_reg_30__8_ ( .D(n2524), .CK(clk_i), .Q(reg_file[40]), .QN(
        n3911) );
  DFF_X1 reg_file_reg_29__8_ ( .D(n2525), .CK(clk_i), .Q(reg_file[72]), .QN(
        n3910) );
  DFF_X1 reg_file_reg_28__8_ ( .D(n2526), .CK(clk_i), .Q(reg_file[104]), .QN(
        n4430) );
  DFF_X1 reg_file_reg_27__8_ ( .D(n2527), .CK(clk_i), .Q(reg_file[136]), .QN(
        n4207) );
  DFF_X1 reg_file_reg_26__8_ ( .D(n2528), .CK(clk_i), .Q(reg_file[168]), .QN(
        n4206) );
  DFF_X1 reg_file_reg_25__8_ ( .D(n2529), .CK(clk_i), .Q(reg_file[200]), .QN(
        n4429) );
  DFF_X1 reg_file_reg_24__8_ ( .D(n2530), .CK(clk_i), .Q(reg_file[232]), .QN(
        n3909) );
  DFF_X1 reg_file_reg_23__8_ ( .D(n2531), .CK(clk_i), .Q(reg_file[264]), .QN(
        n4428) );
  DFF_X1 reg_file_reg_22__8_ ( .D(n2532), .CK(clk_i), .Q(reg_file[296]), .QN(
        n3908) );
  DFF_X1 reg_file_reg_21__8_ ( .D(n2533), .CK(clk_i), .Q(reg_file[328]), .QN(
        n3907) );
  DFF_X1 reg_file_reg_20__8_ ( .D(n2534), .CK(clk_i), .Q(reg_file[360]), .QN(
        n4427) );
  DFF_X1 reg_file_reg_19__8_ ( .D(n2535), .CK(clk_i), .Q(reg_file[392]), .QN(
        n4205) );
  DFF_X1 reg_file_reg_18__8_ ( .D(n2536), .CK(clk_i), .Q(reg_file[424]), .QN(
        n4204) );
  DFF_X1 reg_file_reg_17__8_ ( .D(n2537), .CK(clk_i), .Q(reg_file[456]), .QN(
        n4426) );
  DFF_X1 reg_file_reg_16__8_ ( .D(n2538), .CK(clk_i), .Q(reg_file[488]), .QN(
        n3906) );
  DFF_X1 reg_file_reg_15__8_ ( .D(n2539), .CK(clk_i), .Q(reg_file[520]), .QN(
        n4425) );
  DFF_X1 reg_file_reg_14__8_ ( .D(n2540), .CK(clk_i), .Q(reg_file[552]), .QN(
        n3905) );
  DFF_X1 reg_file_reg_13__8_ ( .D(n2541), .CK(clk_i), .Q(reg_file[584]), .QN(
        n3904) );
  DFF_X1 reg_file_reg_11__8_ ( .D(n2543), .CK(clk_i), .Q(reg_file[648]), .QN(
        n4203) );
  DFF_X1 reg_file_reg_10__8_ ( .D(n2544), .CK(clk_i), .Q(reg_file[680]), .QN(
        n4202) );
  DFF_X1 reg_file_reg_9__8_ ( .D(n2545), .CK(clk_i), .Q(reg_file[712]), .QN(
        n4423) );
  DFF_X1 reg_file_reg_8__8_ ( .D(n2546), .CK(clk_i), .Q(reg_file[744]), .QN(
        n3903) );
  DFF_X1 reg_file_reg_7__8_ ( .D(n2547), .CK(clk_i), .Q(reg_file[776]), .QN(
        n4422) );
  DFF_X1 reg_file_reg_6__8_ ( .D(n2548), .CK(clk_i), .Q(reg_file[808]), .QN(
        n3902) );
  DFF_X1 reg_file_reg_5__8_ ( .D(n2549), .CK(clk_i), .Q(reg_file[840]), .QN(
        n3901) );
  DFF_X1 reg_file_reg_4__8_ ( .D(n2550), .CK(clk_i), .Q(reg_file[872]), .QN(
        n4421) );
  DFF_X1 reg_file_reg_3__8_ ( .D(n2551), .CK(clk_i), .Q(reg_file[904]), .QN(
        n4201) );
  DFF_X1 reg_file_reg_2__8_ ( .D(n2552), .CK(clk_i), .Q(reg_file[936]), .QN(
        n4200) );
  DFF_X1 reg_file_reg_1__8_ ( .D(n2553), .CK(clk_i), .Q(reg_file[968]), .QN(
        n4420) );
  DFF_X1 reg_file_reg_0__8_ ( .D(n2554), .CK(clk_i), .Q(reg_file[1000]), .QN(
        n3900) );
  DFF_X1 reg_file_reg_31__4_ ( .D(n2651), .CK(clk_i), .Q(reg_file[4]) );
  DFF_X1 reg_file_reg_30__4_ ( .D(n2652), .CK(clk_i), .Q(reg_file[36]) );
  DFF_X1 reg_file_reg_29__4_ ( .D(n2653), .CK(clk_i), .Q(reg_file[68]) );
  DFF_X1 reg_file_reg_28__4_ ( .D(n2654), .CK(clk_i), .Q(reg_file[100]) );
  DFF_X1 reg_file_reg_27__4_ ( .D(n2655), .CK(clk_i), .Q(reg_file[132]) );
  DFF_X1 reg_file_reg_26__4_ ( .D(n2656), .CK(clk_i), .Q(reg_file[164]) );
  DFF_X1 reg_file_reg_25__4_ ( .D(n2657), .CK(clk_i), .Q(reg_file[196]) );
  DFF_X1 reg_file_reg_24__4_ ( .D(n2658), .CK(clk_i), .Q(reg_file[228]) );
  DFF_X1 reg_file_reg_23__4_ ( .D(n2659), .CK(clk_i), .Q(reg_file[260]) );
  DFF_X1 reg_file_reg_22__4_ ( .D(n2660), .CK(clk_i), .Q(reg_file[292]) );
  DFF_X1 reg_file_reg_21__4_ ( .D(n2661), .CK(clk_i), .Q(reg_file[324]) );
  DFF_X1 reg_file_reg_20__4_ ( .D(n2662), .CK(clk_i), .Q(reg_file[356]) );
  DFF_X1 reg_file_reg_19__4_ ( .D(n2663), .CK(clk_i), .Q(reg_file[388]) );
  DFF_X1 reg_file_reg_18__4_ ( .D(n2664), .CK(clk_i), .Q(reg_file[420]) );
  DFF_X1 reg_file_reg_17__4_ ( .D(n2665), .CK(clk_i), .Q(reg_file[452]) );
  DFF_X1 reg_file_reg_16__4_ ( .D(n2666), .CK(clk_i), .Q(reg_file[484]) );
  DFF_X1 reg_file_reg_15__4_ ( .D(n2667), .CK(clk_i), .Q(reg_file[516]) );
  DFF_X1 reg_file_reg_14__4_ ( .D(n2668), .CK(clk_i), .Q(reg_file[548]) );
  DFF_X1 reg_file_reg_13__4_ ( .D(n2669), .CK(clk_i), .Q(reg_file[580]) );
  DFF_X1 reg_file_reg_12__4_ ( .D(n2670), .CK(clk_i), .Q(reg_file[612]) );
  DFF_X1 reg_file_reg_11__4_ ( .D(n2671), .CK(clk_i), .Q(reg_file[644]) );
  DFF_X1 reg_file_reg_10__4_ ( .D(n2672), .CK(clk_i), .Q(reg_file[676]) );
  DFF_X1 reg_file_reg_9__4_ ( .D(n2673), .CK(clk_i), .Q(reg_file[708]) );
  DFF_X1 reg_file_reg_8__4_ ( .D(n2674), .CK(clk_i), .Q(reg_file[740]) );
  DFF_X1 reg_file_reg_7__4_ ( .D(n2675), .CK(clk_i), .Q(reg_file[772]) );
  DFF_X1 reg_file_reg_6__4_ ( .D(n2676), .CK(clk_i), .Q(reg_file[804]) );
  DFF_X1 reg_file_reg_5__4_ ( .D(n2677), .CK(clk_i), .Q(reg_file[836]) );
  DFF_X1 reg_file_reg_4__4_ ( .D(n2678), .CK(clk_i), .Q(reg_file[868]) );
  DFF_X1 reg_file_reg_3__4_ ( .D(n2679), .CK(clk_i), .Q(reg_file[900]) );
  DFF_X1 reg_file_reg_2__4_ ( .D(n2680), .CK(clk_i), .Q(reg_file[932]) );
  DFF_X1 reg_file_reg_1__4_ ( .D(n2681), .CK(clk_i), .Q(reg_file[964]) );
  DFF_X1 reg_file_reg_0__4_ ( .D(n2682), .CK(clk_i), .Q(reg_file[996]) );
  DFF_X1 reg_file_reg_31__16_ ( .D(n2267), .CK(clk_i), .Q(reg_file[16]), .QN(
        n4527) );
  DFF_X1 reg_file_reg_30__16_ ( .D(n2268), .CK(clk_i), .Q(reg_file[48]), .QN(
        n4007) );
  DFF_X1 reg_file_reg_29__16_ ( .D(n2269), .CK(clk_i), .Q(reg_file[80]), .QN(
        n4006) );
  DFF_X1 reg_file_reg_28__16_ ( .D(n2270), .CK(clk_i), .Q(reg_file[112]), .QN(
        n4526) );
  DFF_X1 reg_file_reg_27__16_ ( .D(n2271), .CK(clk_i), .Q(reg_file[144]), .QN(
        n4271) );
  DFF_X1 reg_file_reg_26__16_ ( .D(n2272), .CK(clk_i), .Q(reg_file[176]), .QN(
        n4270) );
  DFF_X1 reg_file_reg_25__16_ ( .D(n2273), .CK(clk_i), .Q(reg_file[208]), .QN(
        n4525) );
  DFF_X1 reg_file_reg_24__16_ ( .D(n2274), .CK(clk_i), .Q(reg_file[240]), .QN(
        n4005) );
  DFF_X1 reg_file_reg_23__16_ ( .D(n2275), .CK(clk_i), .Q(reg_file[272]), .QN(
        n4524) );
  DFF_X1 reg_file_reg_22__16_ ( .D(n2276), .CK(clk_i), .Q(reg_file[304]), .QN(
        n4004) );
  DFF_X1 reg_file_reg_21__16_ ( .D(n2277), .CK(clk_i), .Q(reg_file[336]), .QN(
        n4003) );
  DFF_X1 reg_file_reg_20__16_ ( .D(n2278), .CK(clk_i), .Q(reg_file[368]), .QN(
        n4523) );
  DFF_X1 reg_file_reg_19__16_ ( .D(n2279), .CK(clk_i), .Q(reg_file[400]), .QN(
        n4269) );
  DFF_X1 reg_file_reg_18__16_ ( .D(n2280), .CK(clk_i), .Q(reg_file[432]), .QN(
        n4268) );
  DFF_X1 reg_file_reg_17__16_ ( .D(n2281), .CK(clk_i), .Q(reg_file[464]), .QN(
        n4522) );
  DFF_X1 reg_file_reg_16__16_ ( .D(n2282), .CK(clk_i), .Q(reg_file[496]), .QN(
        n4002) );
  DFF_X1 reg_file_reg_15__16_ ( .D(n2283), .CK(clk_i), .Q(reg_file[528]), .QN(
        n4521) );
  DFF_X1 reg_file_reg_14__16_ ( .D(n2284), .CK(clk_i), .Q(reg_file[560]), .QN(
        n4001) );
  DFF_X1 reg_file_reg_13__16_ ( .D(n2285), .CK(clk_i), .Q(reg_file[592]), .QN(
        n4000) );
  DFF_X1 reg_file_reg_12__16_ ( .D(n2286), .CK(clk_i), .Q(reg_file[624]), .QN(
        n4520) );
  DFF_X1 reg_file_reg_11__16_ ( .D(n2287), .CK(clk_i), .Q(reg_file[656]), .QN(
        n4267) );
  DFF_X1 reg_file_reg_10__16_ ( .D(n2288), .CK(clk_i), .Q(reg_file[688]), .QN(
        n4266) );
  DFF_X1 reg_file_reg_9__16_ ( .D(n2289), .CK(clk_i), .Q(reg_file[720]), .QN(
        n4519) );
  DFF_X1 reg_file_reg_8__16_ ( .D(n2290), .CK(clk_i), .Q(reg_file[752]), .QN(
        n3999) );
  DFF_X1 reg_file_reg_7__16_ ( .D(n2291), .CK(clk_i), .Q(reg_file[784]), .QN(
        n4518) );
  DFF_X1 reg_file_reg_6__16_ ( .D(n2292), .CK(clk_i), .Q(reg_file[816]), .QN(
        n3998) );
  DFF_X1 reg_file_reg_5__16_ ( .D(n2293), .CK(clk_i), .Q(reg_file[848]), .QN(
        n3997) );
  DFF_X1 reg_file_reg_4__16_ ( .D(n2294), .CK(clk_i), .Q(reg_file[880]), .QN(
        n4517) );
  DFF_X1 reg_file_reg_3__16_ ( .D(n2295), .CK(clk_i), .Q(reg_file[912]), .QN(
        n4265) );
  DFF_X1 reg_file_reg_2__16_ ( .D(n2296), .CK(clk_i), .Q(reg_file[944]), .QN(
        n4264) );
  DFF_X1 reg_file_reg_1__16_ ( .D(n2297), .CK(clk_i), .Q(reg_file[976]), .QN(
        n4516) );
  DFF_X1 reg_file_reg_0__16_ ( .D(n2298), .CK(clk_i), .Q(reg_file[1008]), .QN(
        n3996) );
  HA_X1 add_x_67_U33 ( .A(rs1_val_gpr_w[0]), .B(u_lsu_N14), .CO(add_x_67_n32), 
        .S(mem_addr_w[0]) );
  FA_X1 add_x_67_U32 ( .A(rs1_val_gpr_w[1]), .B(add_x_67_B_1_), .CI(
        add_x_67_n32), .CO(add_x_67_n31), .S(mem_addr_w[1]) );
  FA_X1 add_x_67_U31 ( .A(rs1_val_gpr_w[2]), .B(u_lsu_N16), .CI(add_x_67_n31), 
        .CO(add_x_67_n30), .S(mem_addr_w[2]) );
  FA_X1 add_x_67_U30 ( .A(add_x_67_n30), .B(add_x_67_B_3_), .CI(n3524), .CO(
        add_x_67_n29), .S(mem_addr_w[3]) );
  FA_X1 add_x_67_U29 ( .A(rs1_val_gpr_w[4]), .B(add_x_67_B_4_), .CI(
        add_x_67_n29), .CO(add_x_67_n28), .S(mem_addr_w[4]) );
  FA_X1 add_x_67_U28 ( .A(rs1_val_gpr_w[5]), .B(mem_i_inst_i[25]), .CI(
        add_x_67_n28), .CO(add_x_67_n27), .S(mem_addr_w[5]) );
  FA_X1 add_x_67_U27 ( .A(rs1_val_gpr_w[6]), .B(mem_i_inst_i[26]), .CI(
        add_x_67_n27), .CO(add_x_67_n26), .S(mem_addr_w[6]) );
  FA_X1 add_x_67_U26 ( .A(n3523), .B(mem_i_inst_i[27]), .CI(add_x_67_n26), 
        .CO(add_x_67_n25), .S(mem_addr_w[7]) );
  FA_X1 add_x_67_U25 ( .A(rs1_val_gpr_w[8]), .B(mem_i_inst_i[28]), .CI(
        add_x_67_n25), .CO(add_x_67_n24), .S(mem_addr_w[8]) );
  FA_X1 add_x_67_U24 ( .A(rs1_val_gpr_w[9]), .B(mem_i_inst_i[29]), .CI(
        add_x_67_n24), .CO(add_x_67_n23), .S(mem_addr_w[9]) );
  FA_X1 add_x_67_U23 ( .A(rs1_val_gpr_w[10]), .B(mem_i_inst_i[30]), .CI(
        add_x_67_n23), .CO(add_x_67_n22), .S(mem_addr_w[10]) );
  FA_X1 add_x_67_U22 ( .A(mem_i_inst_i[31]), .B(rs1_val_gpr_w[11]), .CI(
        add_x_67_n22), .CO(add_x_67_n21), .S(mem_addr_w[11]) );
  FA_X1 add_x_67_U21 ( .A(mem_i_inst_i[31]), .B(rs1_val_gpr_w[12]), .CI(
        add_x_67_n21), .CO(add_x_67_n20), .S(mem_addr_w[12]) );
  FA_X1 add_x_67_U20 ( .A(mem_i_inst_i[31]), .B(rs1_val_gpr_w[13]), .CI(
        add_x_67_n20), .CO(add_x_67_n19), .S(mem_addr_w[13]) );
  FA_X1 add_x_67_U19 ( .A(mem_i_inst_i[31]), .B(rs1_val_gpr_w[14]), .CI(
        add_x_67_n19), .CO(add_x_67_n18), .S(mem_addr_w[14]) );
  FA_X1 add_x_67_U18 ( .A(mem_i_inst_i[31]), .B(rs1_val_gpr_w[15]), .CI(
        add_x_67_n18), .CO(add_x_67_n17), .S(mem_addr_w[15]) );
  FA_X1 add_x_67_U17 ( .A(mem_i_inst_i[31]), .B(rs1_val_gpr_w[16]), .CI(
        add_x_67_n17), .CO(add_x_67_n16), .S(mem_addr_w[16]) );
  FA_X1 add_x_67_U16 ( .A(mem_i_inst_i[31]), .B(rs1_val_gpr_w[17]), .CI(
        add_x_67_n16), .CO(add_x_67_n15), .S(mem_addr_w[17]) );
  FA_X1 add_x_67_U15 ( .A(mem_i_inst_i[31]), .B(rs1_val_gpr_w[18]), .CI(
        add_x_67_n15), .CO(add_x_67_n14), .S(mem_addr_w[18]) );
  FA_X1 add_x_67_U14 ( .A(mem_i_inst_i[31]), .B(rs1_val_gpr_w[19]), .CI(
        add_x_67_n14), .CO(add_x_67_n13), .S(mem_addr_w[19]) );
  FA_X1 add_x_67_U13 ( .A(mem_i_inst_i[31]), .B(rs1_val_gpr_w[20]), .CI(
        add_x_67_n13), .CO(add_x_67_n12), .S(mem_addr_w[20]) );
  FA_X1 add_x_67_U12 ( .A(mem_i_inst_i[31]), .B(rs1_val_gpr_w[21]), .CI(
        add_x_67_n12), .CO(add_x_67_n11), .S(mem_addr_w[21]) );
  FA_X1 add_x_67_U11 ( .A(mem_i_inst_i[31]), .B(rs1_val_gpr_w[22]), .CI(
        add_x_67_n11), .CO(add_x_67_n10), .S(mem_addr_w[22]) );
  FA_X1 add_x_67_U10 ( .A(mem_i_inst_i[31]), .B(rs1_val_gpr_w[23]), .CI(
        add_x_67_n10), .CO(add_x_67_n9), .S(mem_addr_w[23]) );
  FA_X1 add_x_67_U9 ( .A(mem_i_inst_i[31]), .B(rs1_val_gpr_w[24]), .CI(
        add_x_67_n9), .CO(add_x_67_n8), .S(mem_addr_w[24]) );
  FA_X1 add_x_67_U8 ( .A(mem_i_inst_i[31]), .B(rs1_val_gpr_w[25]), .CI(
        add_x_67_n8), .CO(add_x_67_n7), .S(mem_addr_w[25]) );
  FA_X1 add_x_67_U7 ( .A(mem_i_inst_i[31]), .B(rs1_val_gpr_w[26]), .CI(
        add_x_67_n7), .CO(add_x_67_n6), .S(mem_addr_w[26]) );
  FA_X1 add_x_67_U6 ( .A(mem_i_inst_i[31]), .B(rs1_val_gpr_w[27]), .CI(
        add_x_67_n6), .CO(add_x_67_n5), .S(mem_addr_w[27]) );
  FA_X1 add_x_67_U5 ( .A(mem_i_inst_i[31]), .B(rs1_val_gpr_w[28]), .CI(
        add_x_67_n5), .CO(add_x_67_n4), .S(mem_addr_w[28]) );
  FA_X1 add_x_67_U4 ( .A(mem_i_inst_i[31]), .B(rs1_val_gpr_w[29]), .CI(
        add_x_67_n4), .CO(add_x_67_n3), .S(mem_addr_w[29]) );
  FA_X1 add_x_67_U3 ( .A(mem_i_inst_i[31]), .B(rs1_val_gpr_w[30]), .CI(
        add_x_67_n3), .CO(add_x_67_n2), .S(mem_addr_w[30]) );
  XOR2_X1 sub_x_59_U2 ( .A(rs1_val_gpr_w[31]), .B(n3298), .Z(sub_x_59_n1) );
  NOR2_X1 sub_x_59_U18 ( .A1(n3326), .A2(rs1_val_gpr_w[20]), .ZN(sub_x_59_n17)
         );
  NAND2_X1 sub_x_59_U30 ( .A1(n3340), .A2(rs1_val_gpr_w[17]), .ZN(sub_x_59_n29) );
  NOR2_X1 sub_x_59_U29 ( .A1(n3340), .A2(rs1_val_gpr_w[17]), .ZN(sub_x_59_n28)
         );
  NOR2_X1 sub_x_59_U42 ( .A1(n3378), .A2(rs1_val_gpr_w[14]), .ZN(sub_x_59_n41)
         );
  NOR2_X1 sub_x_59_U66 ( .A1(n3382), .A2(rs1_val_gpr_w[8]), .ZN(sub_x_59_n65)
         );
  NAND2_X1 sub_x_59_U78 ( .A1(n3303), .A2(rs1_val_gpr_w[5]), .ZN(sub_x_59_n77)
         );
  NOR2_X1 sub_x_59_U77 ( .A1(n3303), .A2(rs1_val_gpr_w[5]), .ZN(sub_x_59_n76)
         );
  NAND2_X1 sub_x_59_U86 ( .A1(n3299), .A2(rs1_val_gpr_w[3]), .ZN(sub_x_59_n85)
         );
  NOR2_X1 sub_x_59_U95 ( .A1(n3328), .A2(rs1_val_gpr_w[0]), .ZN(sub_x_59_n94)
         );
  NOR2_X1 sub_x_59_U85 ( .A1(n3299), .A2(rs1_val_gpr_w[3]), .ZN(sub_x_59_n84)
         );
  NAND2_X1 sub_x_60_U78 ( .A1(rs2_val_gpr_w[5]), .A2(n3306), .ZN(sub_x_60_n77)
         );
  NOR2_X1 sub_x_60_U77 ( .A1(rs2_val_gpr_w[5]), .A2(n3306), .ZN(sub_x_60_n76)
         );
  NOR2_X1 sub_x_60_U85 ( .A1(rs2_val_gpr_w[3]), .A2(n3288), .ZN(sub_x_60_n84)
         );
  NAND2_X1 sub_x_60_U62 ( .A1(rs2_val_gpr_w[9]), .A2(n3308), .ZN(sub_x_60_n61)
         );
  FA_X1 sub_x_60_U9 ( .A(rs2_val_gpr_w[24]), .B(n3335), .CI(sub_x_60_n9), .CO(
        sub_x_60_n8) );
  FA_X1 DP_OP_181_135_5161_U29 ( .A(DP_OP_181_135_5161_n94), .B(
        DP_OP_181_135_5161_n73), .CI(DP_OP_181_135_5161_n29), .CO(
        DP_OP_181_135_5161_n28), .S(U4_RSOP_173_C3_DATA1_4) );
  FA_X1 DP_OP_181_135_5161_U26 ( .A(DP_OP_181_135_5161_n97), .B(
        DP_OP_181_135_5161_n76), .CI(DP_OP_181_135_5161_n26), .CO(
        DP_OP_181_135_5161_n25), .S(U4_RSOP_173_C3_DATA1_7) );
  FA_X1 DP_OP_181_135_5161_U25 ( .A(DP_OP_181_135_5161_n98), .B(
        DP_OP_181_135_5161_n77), .CI(DP_OP_181_135_5161_n25), .CO(
        DP_OP_181_135_5161_n24), .S(U4_RSOP_173_C3_DATA1_8) );
  FA_X1 DP_OP_181_135_5161_U21 ( .A(DP_OP_181_135_5161_n102), .B(
        DP_OP_181_135_5161_n81), .CI(DP_OP_181_135_5161_n21), .CO(
        DP_OP_181_135_5161_n20), .S(U4_RSOP_173_C3_DATA1_12) );
  FA_X1 DP_OP_181_135_5161_U18 ( .A(DP_OP_181_135_5161_n105), .B(
        DP_OP_181_135_5161_n84), .CI(DP_OP_181_135_5161_n18), .CO(
        DP_OP_181_135_5161_n17), .S(U4_RSOP_173_C3_DATA1_15) );
  FA_X1 DP_OP_181_135_5161_U17 ( .A(DP_OP_181_135_5161_n106), .B(
        DP_OP_181_135_5161_n85), .CI(DP_OP_181_135_5161_n17), .CO(
        DP_OP_181_135_5161_n16), .S(U4_RSOP_173_C3_DATA1_16) );
  FA_X1 DP_OP_181_135_5161_U14 ( .A(DP_OP_181_135_5161_n109), .B(
        DP_OP_181_135_5161_n88), .CI(DP_OP_181_135_5161_n14), .CO(
        DP_OP_181_135_5161_n13), .S(U4_RSOP_173_C3_DATA1_19) );
  FA_X1 DP_OP_181_135_5161_U13 ( .A(DP_OP_181_135_5161_n110), .B(
        DP_OP_181_135_5161_n89), .CI(DP_OP_181_135_5161_n13), .CO(
        DP_OP_181_135_5161_n12), .S(U4_RSOP_173_C3_DATA1_20) );
  FA_X1 DP_OP_181_135_5161_U12 ( .A(DP_OP_181_135_5161_n111), .B(
        DP_OP_181_135_5161_n89), .CI(DP_OP_181_135_5161_n12), .CO(
        DP_OP_181_135_5161_n11), .S(U4_RSOP_173_C3_DATA1_21) );
  FA_X1 DP_OP_181_135_5161_U11 ( .A(DP_OP_181_135_5161_n112), .B(
        DP_OP_181_135_5161_n89), .CI(DP_OP_181_135_5161_n11), .CO(
        DP_OP_181_135_5161_n10), .S(U4_RSOP_173_C3_DATA1_22) );
  FA_X1 DP_OP_181_135_5161_U10 ( .A(DP_OP_181_135_5161_n113), .B(
        DP_OP_181_135_5161_n89), .CI(DP_OP_181_135_5161_n10), .CO(
        DP_OP_181_135_5161_n9), .S(U4_RSOP_173_C3_DATA1_23) );
  FA_X1 DP_OP_181_135_5161_U5 ( .A(DP_OP_181_135_5161_n118), .B(n3391), .CI(
        DP_OP_181_135_5161_n5), .CO(DP_OP_181_135_5161_n4), .S(
        U4_RSOP_173_C3_DATA1_28) );
  FA_X1 DP_OP_181_135_5161_U4 ( .A(DP_OP_181_135_5161_n119), .B(n3391), .CI(
        DP_OP_181_135_5161_n4), .CO(DP_OP_181_135_5161_n3), .S(
        U4_RSOP_173_C3_DATA1_29) );
  OR2_X1 sub_x_60_U29 ( .A1(rs2_val_gpr_w[17]), .A2(n3300), .ZN(sub_x_60_n28)
         );
  AND2_X1 sub_x_60_U30 ( .A1(rs2_val_gpr_w[17]), .A2(n3300), .ZN(sub_x_60_n29)
         );
  OR2_X1 sub_x_60_U13 ( .A1(rs2_val_gpr_w[21]), .A2(n3301), .ZN(sub_x_60_n12)
         );
  DFF_X1 load_signed_q_reg ( .D(n2811), .CK(clk_i), .Q(n3867), .QN(n162) );
  DFF_X1 load_byte_q_reg ( .D(n2815), .CK(clk_i), .Q(n3875), .QN(n158) );
  DFF_X1 alu_func_q_reg_3_ ( .D(n2876), .CK(clk_i), .Q(n3835), .QN(n154) );
  DFF_X1 alu_func_q_reg_1_ ( .D(n2878), .CK(clk_i), .Q(n3765), .QN(n156) );
  DFF_X1 alu_func_q_reg_0_ ( .D(n2879), .CK(clk_i), .Q(n3830), .QN(n157) );
  DFF_X1 alu_func_q_reg_2_ ( .D(n2877), .CK(clk_i), .Q(n3788), .QN(n155) );
  DFF_X1 load_offset_q_reg_0_ ( .D(n2812), .CK(clk_i), .Q(n3874), .QN(n161) );
  DFF_X1 alu_a_q_reg_11_ ( .D(n2799), .CK(clk_i), .Q(alu_a_q[11]), .QN(n3813)
         );
  DFF_X1 alu_a_q_reg_13_ ( .D(n2797), .CK(clk_i), .Q(alu_a_q[13]), .QN(n3815)
         );
  DFF_X1 alu_a_q_reg_15_ ( .D(n2795), .CK(clk_i), .Q(alu_a_q[15]), .QN(n3785)
         );
  DFF_X1 alu_a_q_reg_16_ ( .D(n2794), .CK(clk_i), .Q(alu_a_q[16]), .QN(n3793)
         );
  DFF_X1 alu_a_q_reg_17_ ( .D(n2793), .CK(clk_i), .Q(alu_a_q[17]), .QN(n3794)
         );
  DFF_X1 alu_b_q_reg_28_ ( .D(n2846), .CK(clk_i), .Q(alu_b_q[28]), .QN(n3834)
         );
  DFF_X1 alu_a_q_reg_12_ ( .D(n2798), .CK(clk_i), .Q(alu_a_q[12]), .QN(n3777)
         );
  DFF_X1 alu_a_q_reg_21_ ( .D(n2789), .CK(clk_i), .Q(alu_a_q[21]), .QN(n3766)
         );
  DFF_X1 load_offset_q_reg_1_ ( .D(n2813), .CK(clk_i), .Q(n3866), .QN(n160) );
  DFF_X1 alu_b_q_reg_13_ ( .D(n2861), .CK(clk_i), .Q(alu_b_q[13]), .QN(n3776)
         );
  DFF_X1 alu_b_q_reg_2_ ( .D(n2872), .CK(clk_i), .Q(alu_b_q[2]), .QN(n3763) );
  DFF_X1 alu_b_q_reg_12_ ( .D(n2862), .CK(clk_i), .Q(alu_b_q[12]), .QN(n3806)
         );
  DFF_X1 alu_a_q_reg_19_ ( .D(n2791), .CK(clk_i), .Q(alu_a_q[19]), .QN(n3787)
         );
  DFF_X1 alu_a_q_reg_20_ ( .D(n2790), .CK(clk_i), .Q(alu_a_q[20]), .QN(n3791)
         );
  DFF_X1 alu_a_q_reg_18_ ( .D(n2792), .CK(clk_i), .Q(alu_a_q[18]), .QN(n3786)
         );
  DFF_X1 alu_b_q_reg_10_ ( .D(n2864), .CK(clk_i), .Q(alu_b_q[10]), .QN(n3844)
         );
  DFF_X1 alu_b_q_reg_9_ ( .D(n2865), .CK(clk_i), .Q(alu_b_q[9]), .QN(n3782) );
  DFF_X1 alu_b_q_reg_8_ ( .D(n2866), .CK(clk_i), .Q(alu_b_q[8]), .QN(n3805) );
  DFF_X1 alu_b_q_reg_7_ ( .D(n2867), .CK(clk_i), .Q(alu_b_q[7]), .QN(n3814) );
  DFF_X1 alu_b_q_reg_6_ ( .D(n2868), .CK(clk_i), .Q(alu_b_q[6]), .QN(n3810) );
  DFF_X1 alu_b_q_reg_31_ ( .D(n2843), .CK(clk_i), .Q(alu_b_q[31]), .QN(n3873)
         );
  DFF_X1 alu_b_q_reg_29_ ( .D(n2845), .CK(clk_i), .Q(alu_b_q[29]), .QN(n3836)
         );
  DFF_X1 alu_b_q_reg_27_ ( .D(n2847), .CK(clk_i), .Q(alu_b_q[27]), .QN(n3843)
         );
  DFF_X1 alu_b_q_reg_26_ ( .D(n2848), .CK(clk_i), .Q(alu_b_q[26]), .QN(n3783)
         );
  DFF_X1 alu_b_q_reg_14_ ( .D(n2860), .CK(clk_i), .Q(alu_b_q[14]), .QN(n3846)
         );
  DFF_X1 alu_b_q_reg_11_ ( .D(n2863), .CK(clk_i), .Q(alu_b_q[11]), .QN(n3775)
         );
  DFF_X1 alu_a_q_reg_31_ ( .D(n2779), .CK(clk_i), .Q(alu_a_q[31]), .QN(n3831)
         );
  DFF_X1 alu_a_q_reg_30_ ( .D(n2780), .CK(clk_i), .Q(alu_a_q[30]), .QN(n3833)
         );
  DFF_X1 alu_a_q_reg_29_ ( .D(n2781), .CK(clk_i), .Q(alu_a_q[29]), .QN(n3797)
         );
  DFF_X1 alu_a_q_reg_28_ ( .D(n2782), .CK(clk_i), .Q(alu_a_q[28]), .QN(n3790)
         );
  DFF_X1 alu_a_q_reg_27_ ( .D(n2783), .CK(clk_i), .Q(alu_a_q[27]), .QN(n3784)
         );
  DFF_X1 alu_a_q_reg_26_ ( .D(n2784), .CK(clk_i), .Q(alu_a_q[26]), .QN(n3832)
         );
  DFF_X1 alu_a_q_reg_9_ ( .D(n2801), .CK(clk_i), .Q(alu_a_q[9]), .QN(n3811) );
  DFF_X1 alu_a_q_reg_8_ ( .D(n2802), .CK(clk_i), .Q(alu_a_q[8]), .QN(n3778) );
  DFF_X1 alu_a_q_reg_25_ ( .D(n2785), .CK(clk_i), .Q(alu_a_q[25]), .QN(n3829)
         );
  DFF_X1 alu_a_q_reg_24_ ( .D(n2786), .CK(clk_i), .Q(alu_a_q[24]), .QN(n3789)
         );
  DFF_X1 alu_a_q_reg_23_ ( .D(n2787), .CK(clk_i), .Q(alu_a_q[23]), .QN(n3792)
         );
  DFF_X1 alu_a_q_reg_22_ ( .D(n2788), .CK(clk_i), .Q(alu_a_q[22]), .QN(n3795)
         );
  DFF_X1 alu_a_q_reg_2_ ( .D(n6595), .CK(clk_i), .Q(n3803), .QN(alu_a_q[2]) );
  DFF_X1 alu_a_q_reg_0_ ( .D(n4971), .CK(clk_i), .Q(n3808), .QN(alu_a_q[0]) );
  DFF_X1 alu_a_q_reg_5_ ( .D(n6603), .CK(clk_i), .Q(n3781), .QN(alu_a_q[5]) );
  DFF_X1 alu_a_q_reg_4_ ( .D(n6597), .CK(clk_i), .Q(n3780), .QN(alu_a_q[4]) );
  DFF_X1 alu_a_q_reg_1_ ( .D(n6599), .CK(clk_i), .Q(n3779), .QN(alu_a_q[1]) );
  DFF_X1 alu_a_q_reg_3_ ( .D(n6601), .CK(clk_i), .Q(n3804), .QN(alu_a_q[3]) );
  DFF_X1 alu_b_q_reg_24_ ( .D(n2850), .CK(clk_i), .Q(alu_b_q[24]), .QN(n3840)
         );
  DFF_X1 alu_b_q_reg_23_ ( .D(n2851), .CK(clk_i), .Q(alu_b_q[23]), .QN(n3841)
         );
  DFF_X1 alu_b_q_reg_22_ ( .D(n2852), .CK(clk_i), .Q(alu_b_q[22]), .QN(n3845)
         );
  DFF_X1 alu_b_q_reg_21_ ( .D(n2853), .CK(clk_i), .Q(alu_b_q[21]), .QN(n3839)
         );
  DFF_X1 alu_b_q_reg_20_ ( .D(n2854), .CK(clk_i), .Q(alu_b_q[20]), .QN(n3849)
         );
  DFF_X1 alu_b_q_reg_19_ ( .D(n2855), .CK(clk_i), .Q(alu_b_q[19]), .QN(n3850)
         );
  DFF_X1 alu_b_q_reg_18_ ( .D(n2856), .CK(clk_i), .Q(alu_b_q[18]), .QN(n3838)
         );
  DFF_X1 alu_b_q_reg_17_ ( .D(n2857), .CK(clk_i), .Q(alu_b_q[17]), .QN(n3847)
         );
  DFF_X1 alu_b_q_reg_16_ ( .D(n2858), .CK(clk_i), .Q(alu_b_q[16]), .QN(n3848)
         );
  DFF_X1 alu_b_q_reg_15_ ( .D(n2859), .CK(clk_i), .Q(alu_b_q[15]), .QN(n3851)
         );
  DFF_X1 alu_b_q_reg_4_ ( .D(n2870), .CK(clk_i), .Q(alu_b_q[4]), .QN(n3809) );
  DFF_X1 alu_b_q_reg_5_ ( .D(n2869), .CK(clk_i), .Q(alu_b_q[5]), .QN(n3812) );
  DFF_X1 alu_a_q_reg_6_ ( .D(n2804), .CK(clk_i), .Q(alu_a_q[6]), .QN(n3773) );
  DFF_X1 reg_file_reg_26__7_ ( .D(n2560), .CK(clk_i), .Q(reg_file[167]), .QN(
        n4198) );
  DFF_X1 reg_file_reg_25__7_ ( .D(n2561), .CK(clk_i), .Q(reg_file[199]), .QN(
        n4417) );
  DFF_X1 reg_file_reg_24__7_ ( .D(n2562), .CK(clk_i), .Q(reg_file[231]), .QN(
        n3897) );
  DFF_X1 reg_file_reg_23__7_ ( .D(n2563), .CK(clk_i), .Q(reg_file[263]), .QN(
        n4416) );
  DFF_X1 reg_file_reg_22__7_ ( .D(n2564), .CK(clk_i), .Q(reg_file[295]), .QN(
        n3896) );
  DFF_X1 reg_file_reg_21__7_ ( .D(n2565), .CK(clk_i), .Q(reg_file[327]), .QN(
        n3895) );
  DFF_X1 reg_file_reg_23__6_ ( .D(n2595), .CK(clk_i), .Q(reg_file[262]), .QN(
        n4404) );
  DFF_X1 reg_file_reg_22__6_ ( .D(n2596), .CK(clk_i), .Q(reg_file[294]), .QN(
        n3884) );
  DFF_X1 reg_file_reg_21__6_ ( .D(n2597), .CK(clk_i), .Q(reg_file[326]), .QN(
        n3883) );
  DFF_X1 alu_b_q_reg_3_ ( .D(n6667), .CK(clk_i), .Q(n3772), .QN(alu_b_q[3]) );
  DFF_X1 alu_b_q_reg_1_ ( .D(n6669), .CK(clk_i), .Q(n3807), .QN(alu_b_q[1]) );
  DFF_X1 alu_b_q_reg_0_ ( .D(n6671), .CK(clk_i), .Q(n3774), .QN(alu_b_q[0]) );
  DFF_X1 reg_file_reg_26__6_ ( .D(n2592), .CK(clk_i), .Q(reg_file[166]), .QN(
        n4190) );
  DFF_X1 reg_file_reg_25__6_ ( .D(n2593), .CK(clk_i), .Q(reg_file[198]), .QN(
        n4405) );
  DFF_X1 reg_file_reg_24__6_ ( .D(n2594), .CK(clk_i), .Q(reg_file[230]), .QN(
        n3885) );
  DFF_X1 rd_q_reg_3_ ( .D(n2881), .CK(clk_i), .Q(n3868), .QN(n144) );
  DFF_X1 rd_q_reg_2_ ( .D(n2882), .CK(clk_i), .Q(n3767), .QN(n145) );
  DFF_X1 rd_q_reg_1_ ( .D(n2883), .CK(clk_i), .Q(n3865), .QN(n146) );
  DFF_X1 rd_q_reg_0_ ( .D(n2884), .CK(clk_i), .Q(n3798), .QN(n147) );
  DFF_X1 reg_file_reg_12__8_ ( .D(n2542), .CK(clk_i), .Q(reg_file[616]), .QN(
        n4424) );
  DFF_X1 reg_file_reg_15__7_ ( .D(n2571), .CK(clk_i), .Q(reg_file[519]), .QN(
        n4413) );
  DFF_X1 reg_file_reg_14__7_ ( .D(n2572), .CK(clk_i), .Q(reg_file[551]), .QN(
        n3893) );
  DFF_X1 reg_file_reg_13__7_ ( .D(n2573), .CK(clk_i), .Q(reg_file[583]), .QN(
        n3892) );
  DFF_X1 reg_file_reg_12__7_ ( .D(n2574), .CK(clk_i), .Q(reg_file[615]), .QN(
        n4412) );
  DFF_X1 reg_file_reg_11__7_ ( .D(n2575), .CK(clk_i), .Q(reg_file[647]), .QN(
        n4195) );
  DFF_X1 reg_file_reg_10__7_ ( .D(n2576), .CK(clk_i), .Q(reg_file[679]), .QN(
        n4194) );
  DFF_X1 reg_file_reg_9__7_ ( .D(n2577), .CK(clk_i), .Q(reg_file[711]), .QN(
        n4411) );
  DFF_X1 reg_file_reg_8__7_ ( .D(n2578), .CK(clk_i), .Q(reg_file[743]), .QN(
        n3891) );
  DFF_X1 reg_file_reg_7__7_ ( .D(n2579), .CK(clk_i), .Q(reg_file[775]), .QN(
        n4410) );
  DFF_X1 reg_file_reg_6__7_ ( .D(n2580), .CK(clk_i), .Q(reg_file[807]), .QN(
        n3890) );
  DFF_X1 reg_file_reg_5__7_ ( .D(n2581), .CK(clk_i), .Q(reg_file[839]), .QN(
        n3889) );
  DFF_X1 reg_file_reg_4__7_ ( .D(n2582), .CK(clk_i), .Q(reg_file[871]), .QN(
        n4409) );
  DFF_X1 reg_file_reg_3__7_ ( .D(n2583), .CK(clk_i), .Q(reg_file[903]), .QN(
        n4193) );
  DFF_X1 reg_file_reg_2__7_ ( .D(n2584), .CK(clk_i), .Q(reg_file[935]), .QN(
        n4192) );
  DFF_X1 reg_file_reg_1__7_ ( .D(n2585), .CK(clk_i), .Q(reg_file[967]), .QN(
        n4408) );
  DFF_X1 reg_file_reg_0__7_ ( .D(n2586), .CK(clk_i), .Q(reg_file[999]), .QN(
        n3888) );
  DFF_X1 reg_file_reg_31__7_ ( .D(n2555), .CK(clk_i), .Q(reg_file[7]), .QN(
        n4419) );
  DFF_X1 reg_file_reg_30__7_ ( .D(n2556), .CK(clk_i), .Q(reg_file[39]), .QN(
        n3899) );
  DFF_X1 reg_file_reg_29__7_ ( .D(n2557), .CK(clk_i), .Q(reg_file[71]), .QN(
        n3898) );
  DFF_X1 reg_file_reg_28__7_ ( .D(n2558), .CK(clk_i), .Q(reg_file[103]), .QN(
        n4418) );
  DFF_X1 reg_file_reg_27__7_ ( .D(n2559), .CK(clk_i), .Q(reg_file[135]), .QN(
        n4199) );
  DFF_X1 reg_file_reg_20__7_ ( .D(n2566), .CK(clk_i), .Q(reg_file[359]), .QN(
        n4415) );
  DFF_X1 reg_file_reg_19__7_ ( .D(n2567), .CK(clk_i), .Q(reg_file[391]), .QN(
        n4197) );
  DFF_X1 reg_file_reg_18__7_ ( .D(n2568), .CK(clk_i), .Q(reg_file[423]), .QN(
        n4196) );
  DFF_X1 reg_file_reg_17__7_ ( .D(n2569), .CK(clk_i), .Q(reg_file[455]), .QN(
        n4414) );
  DFF_X1 reg_file_reg_16__7_ ( .D(n2570), .CK(clk_i), .Q(reg_file[487]), .QN(
        n3894) );
  DFF_X1 reg_file_reg_20__6_ ( .D(n2598), .CK(clk_i), .Q(reg_file[358]), .QN(
        n4403) );
  DFF_X1 reg_file_reg_19__6_ ( .D(n2599), .CK(clk_i), .Q(reg_file[390]), .QN(
        n4189) );
  DFF_X1 reg_file_reg_18__6_ ( .D(n2600), .CK(clk_i), .Q(reg_file[422]), .QN(
        n4188) );
  DFF_X1 reg_file_reg_17__6_ ( .D(n2601), .CK(clk_i), .Q(reg_file[454]), .QN(
        n4402) );
  DFF_X1 reg_file_reg_16__6_ ( .D(n2602), .CK(clk_i), .Q(reg_file[486]), .QN(
        n3882) );
  DFF_X1 reg_file_reg_15__6_ ( .D(n2603), .CK(clk_i), .Q(reg_file[518]), .QN(
        n4401) );
  DFF_X1 reg_file_reg_14__6_ ( .D(n2604), .CK(clk_i), .Q(reg_file[550]), .QN(
        n3881) );
  DFF_X1 reg_file_reg_13__6_ ( .D(n2605), .CK(clk_i), .Q(reg_file[582]), .QN(
        n3880) );
  DFF_X1 reg_file_reg_12__6_ ( .D(n2606), .CK(clk_i), .Q(reg_file[614]), .QN(
        n4400) );
  DFF_X1 reg_file_reg_11__6_ ( .D(n2607), .CK(clk_i), .Q(reg_file[646]), .QN(
        n4187) );
  DFF_X1 reg_file_reg_10__6_ ( .D(n2608), .CK(clk_i), .Q(reg_file[678]), .QN(
        n4186) );
  DFF_X1 reg_file_reg_9__6_ ( .D(n2609), .CK(clk_i), .Q(reg_file[710]), .QN(
        n4399) );
  DFF_X1 reg_file_reg_8__6_ ( .D(n2610), .CK(clk_i), .Q(reg_file[742]), .QN(
        n3879) );
  DFF_X1 reg_file_reg_7__6_ ( .D(n2611), .CK(clk_i), .Q(reg_file[774]), .QN(
        n4398) );
  DFF_X1 reg_file_reg_6__6_ ( .D(n2612), .CK(clk_i), .Q(reg_file[806]), .QN(
        n3878) );
  DFF_X1 reg_file_reg_5__6_ ( .D(n2613), .CK(clk_i), .Q(reg_file[838]), .QN(
        n3877) );
  DFF_X1 reg_file_reg_4__6_ ( .D(n2614), .CK(clk_i), .Q(reg_file[870]), .QN(
        n4397) );
  DFF_X1 reg_file_reg_3__6_ ( .D(n2615), .CK(clk_i), .Q(reg_file[902]), .QN(
        n4185) );
  DFF_X1 pc_q_reg_30_ ( .D(n2886), .CK(clk_i), .Q(mem_i_pc_o[30]), .QN(n3870)
         );
  DFF_X1 pc_q_reg_29_ ( .D(n2887), .CK(clk_i), .Q(mem_i_pc_o[29]), .QN(n3871)
         );
  NOR2_X1 U2899 ( .A1(n4945), .A2(mem_i_inst_i[15]), .ZN(n6386) );
  INV_X1 U2900 ( .A(n7774), .ZN(n7743) );
  NAND4_X1 U2901 ( .A1(n5208), .A2(n5209), .A3(n5210), .A4(n5211), .ZN(n2926)
         );
  AOI22_X1 U2902 ( .A1(n3389), .A2(n5207), .B1(n3361), .B2(n2926), .ZN(n2927)
         );
  NAND4_X1 U2903 ( .A1(n5212), .A2(n5213), .A3(n5214), .A4(n5215), .ZN(n2928)
         );
  AOI22_X1 U2904 ( .A1(n3390), .A2(n5220), .B1(n5805), .B2(n2928), .ZN(n2929)
         );
  NAND2_X1 U2905 ( .A1(n2927), .A2(n2929), .ZN(rs2_val_gpr_w[4]) );
  NAND4_X1 U2906 ( .A1(n6229), .A2(n6230), .A3(n6231), .A4(n6232), .ZN(n2930)
         );
  NAND4_X1 U2907 ( .A1(n6233), .A2(n6234), .A3(n6235), .A4(n6236), .ZN(n2931)
         );
  AOI22_X1 U2908 ( .A1(n3387), .A2(n2930), .B1(n3362), .B2(n2931), .ZN(n2932)
         );
  AOI22_X1 U2909 ( .A1(n6373), .A2(n6241), .B1(n3388), .B2(n6246), .ZN(n2933)
         );
  NAND2_X2 U2910 ( .A1(n2932), .A2(n2933), .ZN(rs1_val_gpr_w[19]) );
  AOI22_X1 U2911 ( .A1(reset_vector_i[21]), .A2(n6554), .B1(mem_i_pc_o[21]), 
        .B2(n6588), .ZN(n2934) );
  AOI22_X1 U2912 ( .A1(n3363), .A2(U4_RSOP_173_C3_DATA1_21), .B1(
        csr_mepc_w[21]), .B2(n3319), .ZN(n2935) );
  AOI21_X1 U2913 ( .B1(n6692), .B2(n6693), .A(n6691), .ZN(n2936) );
  NAND2_X1 U2914 ( .A1(n6555), .A2(n2936), .ZN(n2937) );
  NAND3_X1 U2915 ( .A1(n2934), .A2(n2935), .A3(n2937), .ZN(n2895) );
  NOR4_X1 U2916 ( .A1(n3530), .A2(n3612), .A3(n3536), .A4(n3629), .ZN(n2938)
         );
  OAI21_X1 U2917 ( .B1(sub_x_60_n78), .B2(sub_x_60_n76), .A(sub_x_60_n77), 
        .ZN(n2939) );
  NAND2_X1 U2918 ( .A1(n2939), .A2(n2938), .ZN(n3539) );
  AOI22_X1 U2919 ( .A1(n4783), .A2(reg_file[109]), .B1(n4773), .B2(
        reg_file[77]), .ZN(n2940) );
  AOI22_X1 U2920 ( .A1(n3294), .A2(reg_file[173]), .B1(n4764), .B2(
        reg_file[141]), .ZN(n2941) );
  NAND4_X1 U2921 ( .A1(n5425), .A2(n5426), .A3(n2940), .A4(n2941), .ZN(n2942)
         );
  NAND4_X1 U2922 ( .A1(n5427), .A2(n5428), .A3(n5429), .A4(n5430), .ZN(n2943)
         );
  AOI22_X1 U2923 ( .A1(n4754), .A2(n2942), .B1(n3361), .B2(n2943), .ZN(n2944)
         );
  NAND4_X1 U2924 ( .A1(n5435), .A2(n5436), .A3(n5437), .A4(n5438), .ZN(n2945)
         );
  NAND4_X1 U2925 ( .A1(n5431), .A2(n5432), .A3(n5433), .A4(n5434), .ZN(n2946)
         );
  AOI22_X1 U2926 ( .A1(n3390), .A2(n2945), .B1(n3389), .B2(n2946), .ZN(n2947)
         );
  NAND2_X1 U2927 ( .A1(n2944), .A2(n2947), .ZN(rs2_val_gpr_w[13]) );
  NAND4_X1 U2928 ( .A1(n6247), .A2(n6248), .A3(n6249), .A4(n6250), .ZN(n2948)
         );
  AOI22_X1 U2929 ( .A1(n6373), .A2(n2948), .B1(n3388), .B2(n6255), .ZN(n2949)
         );
  AOI22_X1 U2930 ( .A1(n3387), .A2(n6260), .B1(n3362), .B2(n6265), .ZN(n2950)
         );
  NAND2_X2 U2931 ( .A1(n2949), .A2(n2950), .ZN(rs1_val_gpr_w[20]) );
  AOI22_X1 U2932 ( .A1(reset_vector_i[19]), .A2(n6554), .B1(mem_i_pc_o[19]), 
        .B2(n6588), .ZN(n2951) );
  AOI22_X1 U2933 ( .A1(n3363), .A2(U4_RSOP_173_C3_DATA1_19), .B1(
        csr_mepc_w[19]), .B2(n3319), .ZN(n2952) );
  AOI21_X1 U2934 ( .B1(n6695), .B2(n6696), .A(n6694), .ZN(n2953) );
  NAND2_X1 U2935 ( .A1(n6555), .A2(n2953), .ZN(n2954) );
  NAND3_X1 U2936 ( .A1(n2951), .A2(n2952), .A3(n2954), .ZN(n2897) );
  OAI211_X1 U2937 ( .C1(n6459), .C2(n4710), .A(n4709), .B(n4716), .ZN(n6585)
         );
  AOI22_X1 U2938 ( .A1(n4760), .A2(reg_file[229]), .B1(n4756), .B2(
        reg_file[197]), .ZN(n2955) );
  NAND4_X1 U2939 ( .A1(n5253), .A2(n5254), .A3(n2955), .A4(n5255), .ZN(n2956)
         );
  NAND4_X1 U2940 ( .A1(n5256), .A2(n5257), .A3(n5258), .A4(n5259), .ZN(n2957)
         );
  AOI22_X1 U2941 ( .A1(n5805), .A2(n2956), .B1(n3361), .B2(n2957), .ZN(n2958)
         );
  NAND4_X1 U2942 ( .A1(n5264), .A2(n5265), .A3(n5266), .A4(n5267), .ZN(n2959)
         );
  NAND4_X1 U2943 ( .A1(n5260), .A2(n5261), .A3(n5262), .A4(n5263), .ZN(n2960)
         );
  AOI22_X1 U2944 ( .A1(n3390), .A2(n2959), .B1(n3389), .B2(n2960), .ZN(n2961)
         );
  NAND2_X1 U2945 ( .A1(n2958), .A2(n2961), .ZN(rs2_val_gpr_w[5]) );
  AOI22_X1 U2946 ( .A1(n4815), .A2(reg_file[501]), .B1(n4790), .B2(
        reg_file[405]), .ZN(n2962) );
  AOI22_X1 U2947 ( .A1(n3356), .A2(reg_file[469]), .B1(n4795), .B2(
        reg_file[437]), .ZN(n2963) );
  AOI22_X1 U2948 ( .A1(n3359), .A2(reg_file[341]), .B1(n3286), .B2(
        reg_file[373]), .ZN(n2964) );
  AOI22_X1 U2949 ( .A1(n3358), .A2(reg_file[277]), .B1(n4807), .B2(
        reg_file[309]), .ZN(n2965) );
  NAND4_X1 U2950 ( .A1(n2962), .A2(n2963), .A3(n2964), .A4(n2965), .ZN(n2966)
         );
  AOI22_X1 U2951 ( .A1(n3355), .A2(reg_file[661]), .B1(n4815), .B2(
        reg_file[757]), .ZN(n2967) );
  AOI22_X1 U2952 ( .A1(n3356), .A2(reg_file[725]), .B1(n4795), .B2(
        reg_file[693]), .ZN(n2968) );
  AOI22_X1 U2953 ( .A1(n3359), .A2(reg_file[597]), .B1(n3286), .B2(
        reg_file[629]), .ZN(n2969) );
  AOI22_X1 U2954 ( .A1(n3358), .A2(reg_file[533]), .B1(n4809), .B2(
        reg_file[565]), .ZN(n2970) );
  NAND4_X1 U2955 ( .A1(n2967), .A2(n2968), .A3(n2969), .A4(n2970), .ZN(n2971)
         );
  AOI22_X1 U2956 ( .A1(n3387), .A2(n2966), .B1(n3388), .B2(n2971), .ZN(n2972)
         );
  NAND4_X1 U2957 ( .A1(n6266), .A2(n6267), .A3(n6268), .A4(n6269), .ZN(n2973)
         );
  NAND4_X1 U2958 ( .A1(n6270), .A2(n6271), .A3(n6272), .A4(n6273), .ZN(n2974)
         );
  AOI22_X1 U2959 ( .A1(n6373), .A2(n2973), .B1(n3362), .B2(n2974), .ZN(n2975)
         );
  NAND2_X1 U2960 ( .A1(n2972), .A2(n2975), .ZN(rs1_val_gpr_w[21]) );
  AOI22_X1 U2961 ( .A1(reset_vector_i[15]), .A2(n6554), .B1(mem_i_pc_o[15]), 
        .B2(n6588), .ZN(n2976) );
  AOI22_X1 U2962 ( .A1(n3363), .A2(U4_RSOP_173_C3_DATA1_15), .B1(
        csr_mepc_w[15]), .B2(n3319), .ZN(n2977) );
  AOI21_X1 U2963 ( .B1(n6701), .B2(n6702), .A(n6700), .ZN(n2978) );
  NAND2_X1 U2964 ( .A1(n6555), .A2(n2978), .ZN(n2979) );
  NAND3_X1 U2965 ( .A1(n2976), .A2(n2977), .A3(n2979), .ZN(n2901) );
  OAI211_X1 U2966 ( .C1(n3531), .C2(n3612), .A(n3544), .B(sub_x_60_n61), .ZN(
        n2980) );
  NAND2_X1 U2967 ( .A1(sub_x_60_n61), .A2(n3629), .ZN(n2981) );
  NAND3_X1 U2968 ( .A1(n2981), .A2(n2980), .A3(n3535), .ZN(n3538) );
  AND3_X1 U2969 ( .A1(n6686), .A2(n6679), .A3(n6467), .ZN(n6586) );
  NAND4_X1 U2970 ( .A1(n5407), .A2(n5408), .A3(n5409), .A4(n5410), .ZN(n2982)
         );
  NAND4_X1 U2971 ( .A1(n5411), .A2(n5412), .A3(n5413), .A4(n5414), .ZN(n2983)
         );
  AOI22_X1 U2972 ( .A1(n3389), .A2(n2982), .B1(n4754), .B2(n2983), .ZN(n2984)
         );
  AOI22_X1 U2973 ( .A1(n3390), .A2(n5419), .B1(n3361), .B2(n5424), .ZN(n2985)
         );
  NAND2_X1 U2974 ( .A1(n2984), .A2(n2985), .ZN(rs2_val_gpr_w[12]) );
  AOI22_X1 U2975 ( .A1(n3355), .A2(reg_file[662]), .B1(n4815), .B2(
        reg_file[758]), .ZN(n2986) );
  AOI22_X1 U2976 ( .A1(n3356), .A2(reg_file[726]), .B1(n4795), .B2(
        reg_file[694]), .ZN(n2987) );
  AOI22_X1 U2977 ( .A1(n3286), .A2(reg_file[630]), .B1(n3359), .B2(
        reg_file[598]), .ZN(n2988) );
  AOI22_X1 U2978 ( .A1(n4808), .A2(reg_file[566]), .B1(n3358), .B2(
        reg_file[534]), .ZN(n2989) );
  NAND4_X1 U2979 ( .A1(n2986), .A2(n2987), .A3(n2988), .A4(n2989), .ZN(n2990)
         );
  AOI22_X1 U2980 ( .A1(n6396), .A2(reg_file[246]), .B1(n3355), .B2(
        reg_file[150]), .ZN(n2991) );
  AOI22_X1 U2981 ( .A1(n3356), .A2(reg_file[214]), .B1(n4795), .B2(
        reg_file[182]), .ZN(n2992) );
  AOI22_X1 U2982 ( .A1(n3285), .A2(reg_file[118]), .B1(n3359), .B2(
        reg_file[86]), .ZN(n2993) );
  AOI22_X1 U2983 ( .A1(n4807), .A2(reg_file[54]), .B1(n3358), .B2(reg_file[22]), .ZN(n2994) );
  NAND4_X1 U2984 ( .A1(n2991), .A2(n2992), .A3(n2993), .A4(n2994), .ZN(n2995)
         );
  AOI22_X1 U2985 ( .A1(n3388), .A2(n2990), .B1(n6373), .B2(n2995), .ZN(n2996)
         );
  AOI22_X1 U2986 ( .A1(n3355), .A2(reg_file[406]), .B1(n4815), .B2(
        reg_file[502]), .ZN(n2997) );
  AOI22_X1 U2987 ( .A1(n3356), .A2(reg_file[470]), .B1(n4795), .B2(
        reg_file[438]), .ZN(n2998) );
  AOI22_X1 U2988 ( .A1(n3285), .A2(reg_file[374]), .B1(n3359), .B2(
        reg_file[342]), .ZN(n2999) );
  AOI22_X1 U2989 ( .A1(n4809), .A2(reg_file[310]), .B1(n3358), .B2(
        reg_file[278]), .ZN(n3000) );
  NAND4_X1 U2990 ( .A1(n2997), .A2(n2998), .A3(n2999), .A4(n3000), .ZN(n3001)
         );
  AOI22_X1 U2991 ( .A1(n3355), .A2(reg_file[918]), .B1(n3293), .B2(
        reg_file[1014]), .ZN(n3002) );
  AOI22_X1 U2992 ( .A1(n3356), .A2(reg_file[982]), .B1(n4795), .B2(
        reg_file[950]), .ZN(n3003) );
  AOI22_X1 U2993 ( .A1(n3286), .A2(reg_file[886]), .B1(n3359), .B2(
        reg_file[854]), .ZN(n3004) );
  AOI22_X1 U2994 ( .A1(n4809), .A2(reg_file[822]), .B1(n3358), .B2(
        reg_file[790]), .ZN(n3005) );
  NAND4_X1 U2995 ( .A1(n3002), .A2(n3003), .A3(n3004), .A4(n3005), .ZN(n3006)
         );
  AOI22_X1 U2996 ( .A1(n3387), .A2(n3001), .B1(n3362), .B2(n3006), .ZN(n3007)
         );
  NAND2_X1 U2997 ( .A1(n2996), .A2(n3007), .ZN(rs1_val_gpr_w[22]) );
  AOI22_X1 U2998 ( .A1(reset_vector_i[11]), .A2(n6554), .B1(mem_i_pc_o[11]), 
        .B2(n6588), .ZN(n3008) );
  AOI22_X1 U2999 ( .A1(n3363), .A2(U4_RSOP_173_C3_DATA1_11), .B1(
        csr_mepc_w[11]), .B2(n6589), .ZN(n3009) );
  AOI21_X1 U3000 ( .B1(n6707), .B2(n6708), .A(n6706), .ZN(n3010) );
  NAND2_X1 U3001 ( .A1(n6555), .A2(n3010), .ZN(n3011) );
  NAND3_X1 U3002 ( .A1(n3008), .A2(n3009), .A3(n3011), .ZN(n2905) );
  AOI22_X1 U3003 ( .A1(n4755), .A2(reg_file[463]), .B1(n4758), .B2(
        reg_file[495]), .ZN(n3012) );
  AOI22_X1 U3004 ( .A1(n3294), .A2(reg_file[431]), .B1(n4765), .B2(
        reg_file[399]), .ZN(n3013) );
  AOI22_X1 U3005 ( .A1(n4774), .A2(reg_file[335]), .B1(n5811), .B2(
        reg_file[367]), .ZN(n3014) );
  AOI22_X1 U3006 ( .A1(n4787), .A2(reg_file[303]), .B1(n3296), .B2(
        reg_file[271]), .ZN(n3015) );
  NAND4_X1 U3007 ( .A1(n3012), .A2(n3013), .A3(n3014), .A4(n3015), .ZN(n3016)
         );
  NAND4_X1 U3008 ( .A1(n5456), .A2(n5457), .A3(n5458), .A4(n5459), .ZN(n3017)
         );
  AOI22_X1 U3009 ( .A1(n3389), .A2(n3016), .B1(n4754), .B2(n3017), .ZN(n3018)
         );
  NAND4_X1 U3010 ( .A1(n5460), .A2(n5461), .A3(n5462), .A4(n5463), .ZN(n3019)
         );
  NAND4_X1 U3011 ( .A1(n5464), .A2(n5465), .A3(n5466), .A4(n5467), .ZN(n3020)
         );
  AOI22_X1 U3012 ( .A1(n3390), .A2(n3019), .B1(n3361), .B2(n3020), .ZN(n3021)
         );
  NAND2_X1 U3013 ( .A1(n3018), .A2(n3021), .ZN(rs2_val_gpr_w[15]) );
  AOI22_X1 U3014 ( .A1(n3355), .A2(reg_file[408]), .B1(n3293), .B2(
        reg_file[504]), .ZN(n3022) );
  AOI22_X1 U3015 ( .A1(n3360), .A2(reg_file[440]), .B1(n4800), .B2(
        reg_file[472]), .ZN(n3023) );
  AOI22_X1 U3016 ( .A1(n3285), .A2(reg_file[376]), .B1(n4805), .B2(
        reg_file[344]), .ZN(n3024) );
  AOI22_X1 U3017 ( .A1(n4808), .A2(reg_file[312]), .B1(n4812), .B2(
        reg_file[280]), .ZN(n3025) );
  NAND4_X1 U3018 ( .A1(n3022), .A2(n3023), .A3(n3024), .A4(n3025), .ZN(n3026)
         );
  AOI22_X1 U3019 ( .A1(n4813), .A2(reg_file[1016]), .B1(n3355), .B2(
        reg_file[920]), .ZN(n3027) );
  AOI22_X1 U3020 ( .A1(n3360), .A2(reg_file[952]), .B1(n4800), .B2(
        reg_file[984]), .ZN(n3028) );
  AOI22_X1 U3021 ( .A1(n3286), .A2(reg_file[888]), .B1(n4805), .B2(
        reg_file[856]), .ZN(n3029) );
  AOI22_X1 U3022 ( .A1(n4807), .A2(reg_file[824]), .B1(n4811), .B2(
        reg_file[792]), .ZN(n3030) );
  NAND4_X1 U3023 ( .A1(n3027), .A2(n3028), .A3(n3029), .A4(n3030), .ZN(n3031)
         );
  AOI22_X1 U3024 ( .A1(n3387), .A2(n3026), .B1(n3362), .B2(n3031), .ZN(n3032)
         );
  AOI22_X1 U3025 ( .A1(n3386), .A2(reg_file[664]), .B1(n3293), .B2(
        reg_file[760]), .ZN(n3033) );
  AOI22_X1 U3026 ( .A1(n3360), .A2(reg_file[696]), .B1(n4800), .B2(
        reg_file[728]), .ZN(n3034) );
  AOI22_X1 U3027 ( .A1(n3285), .A2(reg_file[632]), .B1(n4805), .B2(
        reg_file[600]), .ZN(n3035) );
  AOI22_X1 U3028 ( .A1(n4808), .A2(reg_file[568]), .B1(n4811), .B2(
        reg_file[536]), .ZN(n3036) );
  NAND4_X1 U3029 ( .A1(n3033), .A2(n3034), .A3(n3035), .A4(n3036), .ZN(n3037)
         );
  AOI22_X1 U3030 ( .A1(n3355), .A2(reg_file[152]), .B1(n4814), .B2(
        reg_file[248]), .ZN(n3038) );
  AOI22_X1 U3031 ( .A1(n3360), .A2(reg_file[184]), .B1(n4800), .B2(
        reg_file[216]), .ZN(n3039) );
  AOI22_X1 U3032 ( .A1(n3286), .A2(reg_file[120]), .B1(n4805), .B2(
        reg_file[88]), .ZN(n3040) );
  AOI22_X1 U3033 ( .A1(n4807), .A2(reg_file[56]), .B1(n4812), .B2(reg_file[24]), .ZN(n3041) );
  NAND4_X1 U3034 ( .A1(n3038), .A2(n3039), .A3(n3040), .A4(n3041), .ZN(n3042)
         );
  AOI22_X1 U3035 ( .A1(n3388), .A2(n3037), .B1(n6373), .B2(n3042), .ZN(n3043)
         );
  NAND2_X1 U3036 ( .A1(n3032), .A2(n3043), .ZN(rs1_val_gpr_w[24]) );
  INV_X1 U3037 ( .A(reset_vector_i[10]), .ZN(n3044) );
  INV_X1 U3038 ( .A(n6709), .ZN(n3045) );
  AOI221_X1 U3039 ( .B1(reset_vector_i[10]), .B2(n6709), .C1(n3044), .C2(n3045), .A(n6551), .ZN(n3046) );
  AOI21_X1 U3040 ( .B1(n3319), .B2(csr_mepc_w[10]), .A(n3046), .ZN(n3047) );
  AOI22_X1 U3041 ( .A1(reset_vector_i[10]), .A2(n6554), .B1(mem_i_pc_o[10]), 
        .B2(n6588), .ZN(n3048) );
  INV_X1 U3042 ( .A(n3395), .ZN(n3049) );
  AOI21_X1 U3043 ( .B1(n3424), .B2(DP_OP_181_135_5161_n24), .A(n3049), .ZN(
        n3050) );
  XNOR2_X1 U3044 ( .A(DP_OP_181_135_5161_n100), .B(n3050), .ZN(n3051) );
  NAND2_X1 U3045 ( .A1(DP_OP_181_135_5161_n79), .A2(n3051), .ZN(n3052) );
  OAI211_X1 U3046 ( .C1(DP_OP_181_135_5161_n79), .C2(n3051), .A(n3363), .B(
        n3052), .ZN(n3053) );
  NAND3_X1 U3047 ( .A1(n3047), .A2(n3048), .A3(n3053), .ZN(n2906) );
  OAI211_X1 U3048 ( .C1(n6459), .C2(n4710), .A(n4709), .B(n6458), .ZN(n6465)
         );
  NAND4_X1 U3049 ( .A1(n5439), .A2(n5440), .A3(n5441), .A4(n5442), .ZN(n3054)
         );
  NAND4_X1 U3050 ( .A1(n5443), .A2(n5444), .A3(n5445), .A4(n5446), .ZN(n3055)
         );
  AOI22_X1 U3051 ( .A1(n4754), .A2(n3054), .B1(n3361), .B2(n3055), .ZN(n3056)
         );
  NAND4_X1 U3052 ( .A1(n5447), .A2(n5448), .A3(n5449), .A4(n5450), .ZN(n3057)
         );
  AOI22_X1 U3053 ( .A1(n3390), .A2(n5455), .B1(n3389), .B2(n3057), .ZN(n3058)
         );
  NAND2_X2 U3054 ( .A1(n3056), .A2(n3058), .ZN(rs2_val_gpr_w[14]) );
  AOI22_X1 U3055 ( .A1(n4809), .A2(reg_file[313]), .B1(n4811), .B2(
        reg_file[281]), .ZN(n3059) );
  NAND4_X1 U3056 ( .A1(n6298), .A2(n6299), .A3(n3059), .A4(n6300), .ZN(n3060)
         );
  AOI22_X1 U3057 ( .A1(n3355), .A2(reg_file[153]), .B1(n4814), .B2(
        reg_file[249]), .ZN(n3061) );
  AOI22_X1 U3058 ( .A1(n4800), .A2(reg_file[217]), .B1(n3360), .B2(
        reg_file[185]), .ZN(n3062) );
  AOI22_X1 U3059 ( .A1(n3286), .A2(reg_file[121]), .B1(n4805), .B2(
        reg_file[89]), .ZN(n3063) );
  AOI22_X1 U3060 ( .A1(n4812), .A2(reg_file[25]), .B1(n4809), .B2(reg_file[57]), .ZN(n3064) );
  NAND4_X1 U3061 ( .A1(n3061), .A2(n3062), .A3(n3063), .A4(n3064), .ZN(n3065)
         );
  AOI22_X1 U3062 ( .A1(n3387), .A2(n3060), .B1(n6373), .B2(n3065), .ZN(n3066)
         );
  NAND4_X1 U3063 ( .A1(n6301), .A2(n6302), .A3(n6303), .A4(n6304), .ZN(n3067)
         );
  NAND4_X1 U3064 ( .A1(n6305), .A2(n6306), .A3(n6307), .A4(n6308), .ZN(n3068)
         );
  AOI22_X1 U3065 ( .A1(n3388), .A2(n3067), .B1(n3362), .B2(n3068), .ZN(n3069)
         );
  NAND2_X1 U3066 ( .A1(n3066), .A2(n3069), .ZN(rs1_val_gpr_w[25]) );
  AOI22_X1 U3067 ( .A1(reset_vector_i[9]), .A2(n6554), .B1(mem_i_pc_o[9]), 
        .B2(n6588), .ZN(n3070) );
  AOI21_X1 U3068 ( .B1(n6710), .B2(n6711), .A(n6709), .ZN(n3071) );
  AOI22_X1 U3069 ( .A1(n6555), .A2(n3071), .B1(csr_mepc_w[9]), .B2(n6589), 
        .ZN(n3072) );
  XOR2_X1 U3070 ( .A(DP_OP_181_135_5161_n99), .B(DP_OP_181_135_5161_n78), .Z(
        n3073) );
  NAND2_X1 U3071 ( .A1(DP_OP_181_135_5161_n24), .A2(n3073), .ZN(n3074) );
  OAI211_X1 U3072 ( .C1(DP_OP_181_135_5161_n24), .C2(n3073), .A(n3363), .B(
        n3074), .ZN(n3075) );
  NAND3_X1 U3073 ( .A1(n3070), .A2(n3072), .A3(n3075), .ZN(n2907) );
  OAI21_X1 U3074 ( .B1(rs1_val_gpr_w[18]), .B2(n3337), .A(n3594), .ZN(n3076)
         );
  NOR2_X1 U3075 ( .A1(sub_x_59_n17), .A2(n3076), .ZN(n3077) );
  NAND2_X1 U3076 ( .A1(n3595), .A2(n3077), .ZN(n3512) );
  AND3_X1 U3077 ( .A1(n3351), .A2(n3557), .A3(rs2_val_gpr_w[12]), .ZN(n3078)
         );
  AOI21_X1 U3078 ( .B1(n3290), .B2(rs2_val_gpr_w[13]), .A(n3078), .ZN(n3079)
         );
  NAND2_X1 U3079 ( .A1(n3323), .A2(rs2_val_gpr_w[14]), .ZN(n3080) );
  OAI21_X1 U3080 ( .B1(n3079), .B2(n3554), .A(n3080), .ZN(n3529) );
  NAND4_X1 U3081 ( .A1(n5364), .A2(n5365), .A3(n5366), .A4(n5367), .ZN(n3081)
         );
  AOI22_X1 U3082 ( .A1(n5805), .A2(n3081), .B1(n3361), .B2(n5372), .ZN(n3082)
         );
  AOI22_X1 U3083 ( .A1(n3389), .A2(n5377), .B1(n3390), .B2(n5382), .ZN(n3083)
         );
  NAND2_X2 U3084 ( .A1(n3082), .A2(n3083), .ZN(rs2_val_gpr_w[10]) );
  XNOR2_X1 U3085 ( .A(DP_OP_181_135_5161_n121), .B(DP_OP_181_135_5161_n89), 
        .ZN(n3084) );
  NAND2_X1 U3086 ( .A1(n3483), .A2(n3084), .ZN(n3085) );
  OAI211_X1 U3087 ( .C1(n3483), .C2(n3084), .A(n3363), .B(n3085), .ZN(n3454)
         );
  OAI22_X1 U3088 ( .A1(n3289), .A2(n3297), .B1(n4819), .B2(n3820), .ZN(n3086)
         );
  OAI21_X1 U3089 ( .B1(n6585), .B2(n7986), .A(n6562), .ZN(n3087) );
  OAI21_X1 U3090 ( .B1(n3087), .B2(n3086), .A(DP_OP_181_135_5161_n22), .ZN(
        n3088) );
  NAND2_X1 U3091 ( .A1(n3087), .A2(n3086), .ZN(n3089) );
  NAND2_X1 U3092 ( .A1(n3088), .A2(n3089), .ZN(DP_OP_181_135_5161_n21) );
  XNOR2_X1 U3093 ( .A(DP_OP_181_135_5161_n22), .B(n3087), .ZN(n3090) );
  XNOR2_X1 U3094 ( .A(n3090), .B(n3086), .ZN(U4_RSOP_173_C3_DATA1_11) );
  AOI22_X1 U3095 ( .A1(n3293), .A2(reg_file[763]), .B1(n4790), .B2(
        reg_file[667]), .ZN(n3091) );
  AOI22_X1 U3096 ( .A1(n4801), .A2(reg_file[731]), .B1(n4796), .B2(
        reg_file[699]), .ZN(n3092) );
  AOI22_X1 U3097 ( .A1(n3286), .A2(reg_file[635]), .B1(n4806), .B2(
        reg_file[603]), .ZN(n3093) );
  AOI22_X1 U3098 ( .A1(n4811), .A2(reg_file[539]), .B1(n4809), .B2(
        reg_file[571]), .ZN(n3094) );
  NAND4_X1 U3099 ( .A1(n3091), .A2(n3092), .A3(n3093), .A4(n3094), .ZN(n3095)
         );
  NAND4_X1 U3100 ( .A1(n6333), .A2(n6334), .A3(n6335), .A4(n6336), .ZN(n3096)
         );
  AOI22_X1 U3101 ( .A1(n3388), .A2(n3095), .B1(n3362), .B2(n3096), .ZN(n3097)
         );
  AOI22_X1 U3102 ( .A1(n4809), .A2(reg_file[315]), .B1(n4812), .B2(
        reg_file[283]), .ZN(n3098) );
  AOI22_X1 U3103 ( .A1(n4806), .A2(reg_file[347]), .B1(n3285), .B2(
        reg_file[379]), .ZN(n3099) );
  NAND4_X1 U3104 ( .A1(n6337), .A2(n6338), .A3(n3098), .A4(n3099), .ZN(n3100)
         );
  AOI22_X1 U3105 ( .A1(n3355), .A2(reg_file[155]), .B1(n4814), .B2(
        reg_file[251]), .ZN(n3101) );
  AOI22_X1 U3106 ( .A1(n4801), .A2(reg_file[219]), .B1(n4796), .B2(
        reg_file[187]), .ZN(n3102) );
  AOI22_X1 U3107 ( .A1(n4806), .A2(reg_file[91]), .B1(n3285), .B2(
        reg_file[123]), .ZN(n3103) );
  AOI22_X1 U3108 ( .A1(n4809), .A2(reg_file[59]), .B1(n4812), .B2(reg_file[27]), .ZN(n3104) );
  NAND4_X1 U3109 ( .A1(n3101), .A2(n3102), .A3(n3103), .A4(n3104), .ZN(n3105)
         );
  AOI22_X1 U3110 ( .A1(n3387), .A2(n3100), .B1(n6373), .B2(n3105), .ZN(n3106)
         );
  NAND2_X1 U3111 ( .A1(n3097), .A2(n3106), .ZN(rs1_val_gpr_w[27]) );
  AOI22_X1 U3112 ( .A1(reset_vector_i[7]), .A2(n6554), .B1(mem_i_pc_o[7]), 
        .B2(n6588), .ZN(n3107) );
  AOI22_X1 U3113 ( .A1(n3363), .A2(U4_RSOP_173_C3_DATA1_7), .B1(csr_mepc_w[7]), 
        .B2(n6589), .ZN(n3108) );
  AOI21_X1 U3114 ( .B1(n6713), .B2(n6714), .A(n6712), .ZN(n3109) );
  NAND2_X1 U3115 ( .A1(n6555), .A2(n3109), .ZN(n3110) );
  NAND3_X1 U3116 ( .A1(n3107), .A2(n3108), .A3(n3110), .ZN(n2909) );
  OAI211_X1 U3117 ( .C1(rs1_val_gpr_w[10]), .C2(n3381), .A(n3599), .B(n3593), 
        .ZN(n3111) );
  INV_X1 U3118 ( .A(n3111), .ZN(n3583) );
  AND3_X1 U3119 ( .A1(rs1_val_gpr_w[18]), .A2(n3594), .A3(n3337), .ZN(n3112)
         );
  AOI21_X1 U3120 ( .B1(rs1_val_gpr_w[19]), .B2(n3332), .A(n3112), .ZN(n3113)
         );
  NAND2_X1 U3121 ( .A1(rs1_val_gpr_w[20]), .A2(n3326), .ZN(n3114) );
  OAI21_X1 U3122 ( .B1(n3113), .B2(sub_x_59_n17), .A(n3114), .ZN(n3572) );
  NAND3_X1 U3123 ( .A1(n3538), .A2(n3539), .A3(n3537), .ZN(n3115) );
  NAND3_X1 U3124 ( .A1(n3528), .A2(n3555), .A3(n3115), .ZN(n3116) );
  AOI21_X1 U3125 ( .B1(n3555), .B2(n3529), .A(n3545), .ZN(n3117) );
  NAND2_X1 U3126 ( .A1(n3116), .A2(n3117), .ZN(n3527) );
  NAND2_X1 U3127 ( .A1(n3376), .A2(rs1_val_gpr_w[27]), .ZN(n3118) );
  NAND3_X1 U3128 ( .A1(rs1_val_gpr_w[26]), .A2(n3385), .A3(n3488), .ZN(n3119)
         );
  NAND2_X1 U3129 ( .A1(n3119), .A2(n3118), .ZN(n3120) );
  AOI22_X1 U3130 ( .A1(n3348), .A2(rs1_val_gpr_w[28]), .B1(n3477), .B2(n3120), 
        .ZN(n3413) );
  INV_X1 U3131 ( .A(n6586), .ZN(n3121) );
  OAI21_X1 U3132 ( .B1(n6466), .B2(n6579), .A(mem_i_pc_o[1]), .ZN(n3122) );
  OAI21_X1 U3133 ( .B1(n3380), .B2(n3121), .A(n3122), .ZN(
        DP_OP_181_135_5161_n91) );
  AOI22_X1 U3134 ( .A1(n4809), .A2(reg_file[319]), .B1(n4811), .B2(
        reg_file[287]), .ZN(n3123) );
  NAND4_X1 U3135 ( .A1(n6378), .A2(n6379), .A3(n3123), .A4(n6380), .ZN(n3124)
         );
  NAND4_X1 U3136 ( .A1(n6388), .A2(n6389), .A3(n6390), .A4(n6391), .ZN(n3125)
         );
  AOI22_X1 U3137 ( .A1(n3387), .A2(n3124), .B1(n3388), .B2(n3125), .ZN(n3126)
         );
  NAND4_X1 U3138 ( .A1(n6369), .A2(n6370), .A3(n6371), .A4(n6372), .ZN(n3127)
         );
  NAND4_X1 U3139 ( .A1(n6374), .A2(n6375), .A3(n6376), .A4(n6377), .ZN(n3128)
         );
  AOI22_X1 U3140 ( .A1(n6373), .A2(n3127), .B1(n3362), .B2(n3128), .ZN(n3129)
         );
  NAND2_X1 U3141 ( .A1(n3126), .A2(n3129), .ZN(rs1_val_gpr_w[31]) );
  NOR2_X1 U3142 ( .A1(n_0_net__4_), .A2(n6715), .ZN(n3130) );
  OAI21_X1 U3143 ( .B1(reset_vector_i[6]), .B2(n3130), .A(n6714), .ZN(n3131)
         );
  AOI22_X1 U3144 ( .A1(n3319), .A2(csr_mepc_w[6]), .B1(n6588), .B2(
        mem_i_pc_o[6]), .ZN(n3132) );
  XOR2_X1 U3145 ( .A(n3457), .B(DP_OP_181_135_5161_n96), .Z(n3133) );
  XNOR2_X1 U3146 ( .A(n3133), .B(DP_OP_181_135_5161_n75), .ZN(n3134) );
  AOI22_X1 U3147 ( .A1(reset_vector_i[6]), .A2(n6554), .B1(n6559), .B2(n3134), 
        .ZN(n3135) );
  OAI211_X1 U3148 ( .C1(n6551), .C2(n3131), .A(n3132), .B(n3135), .ZN(n2910)
         );
  OAI21_X1 U3149 ( .B1(rs2_val_gpr_w[12]), .B2(n3351), .A(n3557), .ZN(n3136)
         );
  NOR2_X1 U3150 ( .A1(n3554), .A2(n3136), .ZN(n3528) );
  OAI211_X1 U3151 ( .C1(n3339), .C2(rs2_val_gpr_w[16]), .A(n3550), .B(
        sub_x_60_n28), .ZN(n3137) );
  NOR3_X1 U3152 ( .A1(n3648), .A2(n3549), .A3(n3137), .ZN(n3503) );
  OAI21_X1 U3153 ( .B1(n3333), .B2(rs2_val_gpr_w[26]), .A(n3481), .ZN(n3138)
         );
  NOR2_X1 U3154 ( .A1(n3662), .A2(n3138), .ZN(n3416) );
  AOI22_X1 U3155 ( .A1(n4815), .A2(reg_file[751]), .B1(n3386), .B2(
        reg_file[655]), .ZN(n3139) );
  AOI22_X1 U3156 ( .A1(n3314), .A2(reg_file[719]), .B1(n4794), .B2(
        reg_file[687]), .ZN(n3140) );
  AOI22_X1 U3157 ( .A1(n3286), .A2(reg_file[623]), .B1(n3359), .B2(
        reg_file[591]), .ZN(n3141) );
  AOI22_X1 U3158 ( .A1(n3316), .A2(reg_file[527]), .B1(n3315), .B2(
        reg_file[559]), .ZN(n3142) );
  NAND4_X1 U3159 ( .A1(n3139), .A2(n3140), .A3(n3141), .A4(n3142), .ZN(n3143)
         );
  AOI22_X1 U3160 ( .A1(n3316), .A2(reg_file[783]), .B1(n3315), .B2(
        reg_file[815]), .ZN(n3144) );
  AOI22_X1 U3161 ( .A1(n3359), .A2(reg_file[847]), .B1(n3285), .B2(
        reg_file[879]), .ZN(n3145) );
  NAND4_X1 U3162 ( .A1(n6147), .A2(n6148), .A3(n3144), .A4(n3145), .ZN(n3146)
         );
  AOI22_X1 U3163 ( .A1(n3388), .A2(n3143), .B1(n3362), .B2(n3146), .ZN(n3147)
         );
  NAND4_X1 U3164 ( .A1(n6149), .A2(n6150), .A3(n6151), .A4(n6152), .ZN(n3148)
         );
  NAND4_X1 U3165 ( .A1(n6153), .A2(n6154), .A3(n6155), .A4(n6156), .ZN(n3149)
         );
  AOI22_X1 U3166 ( .A1(n6373), .A2(n3148), .B1(n3387), .B2(n3149), .ZN(n3150)
         );
  NAND2_X1 U3167 ( .A1(n3147), .A2(n3150), .ZN(rs1_val_gpr_w[15]) );
  AOI22_X1 U3168 ( .A1(n5809), .A2(reg_file[479]), .B1(n4758), .B2(
        reg_file[511]), .ZN(n3151) );
  AOI22_X1 U3169 ( .A1(n4818), .A2(reg_file[447]), .B1(n3769), .B2(
        reg_file[415]), .ZN(n3152) );
  AOI22_X1 U3170 ( .A1(n4778), .A2(reg_file[383]), .B1(n3799), .B2(
        reg_file[351]), .ZN(n3153) );
  AOI22_X1 U3171 ( .A1(n4788), .A2(reg_file[287]), .B1(n4787), .B2(
        reg_file[319]), .ZN(n3154) );
  NAND4_X1 U3172 ( .A1(n3151), .A2(n3152), .A3(n3153), .A4(n3154), .ZN(n3155)
         );
  AOI22_X1 U3173 ( .A1(n4758), .A2(reg_file[255]), .B1(n4756), .B2(
        reg_file[223]), .ZN(n3156) );
  AOI22_X1 U3174 ( .A1(n4818), .A2(reg_file[191]), .B1(n3769), .B2(
        reg_file[159]), .ZN(n3157) );
  AOI22_X1 U3175 ( .A1(n4778), .A2(reg_file[127]), .B1(n3799), .B2(
        reg_file[95]), .ZN(n3158) );
  AOI22_X1 U3176 ( .A1(n4788), .A2(reg_file[31]), .B1(n4787), .B2(reg_file[63]), .ZN(n3159) );
  NAND4_X1 U3177 ( .A1(n3156), .A2(n3157), .A3(n3158), .A4(n3159), .ZN(n3160)
         );
  AOI22_X1 U3178 ( .A1(n5804), .A2(n3155), .B1(n5805), .B2(n3160), .ZN(n3161)
         );
  AOI22_X1 U3179 ( .A1(n4758), .A2(reg_file[767]), .B1(n3519), .B2(
        reg_file[735]), .ZN(n3162) );
  AOI22_X1 U3180 ( .A1(n4788), .A2(reg_file[543]), .B1(n4787), .B2(
        reg_file[575]), .ZN(n3163) );
  NAND4_X1 U3181 ( .A1(n5807), .A2(n5806), .A3(n3162), .A4(n3163), .ZN(n3164)
         );
  NAND3_X1 U3182 ( .A1(n5814), .A2(n3411), .A3(n5817), .ZN(n3165) );
  AOI22_X1 U3183 ( .A1(n5808), .A2(n3164), .B1(n4816), .B2(n3165), .ZN(n3166)
         );
  NAND2_X1 U3184 ( .A1(n3161), .A2(n3166), .ZN(rs2_val_gpr_w[31]) );
  NOR2_X1 U3185 ( .A1(n3297), .A2(n3526), .ZN(n3167) );
  NOR3_X1 U3186 ( .A1(n6465), .A2(n3801), .A3(n6464), .ZN(n3168) );
  AOI211_X1 U3187 ( .C1(mem_i_pc_o[0]), .C2(n6466), .A(n3167), .B(n3168), .ZN(
        n3169) );
  NOR3_X1 U3188 ( .A1(n6623), .A2(n3297), .A3(n3169), .ZN(
        DP_OP_181_135_5161_n32) );
  NOR2_X1 U3189 ( .A1(n6623), .A2(n3297), .ZN(n3170) );
  XNOR2_X1 U3190 ( .A(n3169), .B(n3170), .ZN(U4_RSOP_173_C3_DATA1_0) );
  AOI22_X1 U3191 ( .A1(n3355), .A2(reg_file[670]), .B1(n4814), .B2(
        reg_file[766]), .ZN(n3171) );
  AOI22_X1 U3192 ( .A1(n4801), .A2(reg_file[734]), .B1(n4797), .B2(
        reg_file[702]), .ZN(n3172) );
  AOI22_X1 U3193 ( .A1(n3286), .A2(reg_file[638]), .B1(n4806), .B2(
        reg_file[606]), .ZN(n3173) );
  AOI22_X1 U3194 ( .A1(n4811), .A2(reg_file[542]), .B1(n4809), .B2(
        reg_file[574]), .ZN(n3174) );
  NAND4_X1 U3195 ( .A1(n3171), .A2(n3172), .A3(n3173), .A4(n3174), .ZN(n3175)
         );
  AOI22_X1 U3196 ( .A1(n4809), .A2(reg_file[62]), .B1(n4812), .B2(reg_file[30]), .ZN(n3176) );
  AOI22_X1 U3197 ( .A1(n3286), .A2(reg_file[126]), .B1(n4806), .B2(
        reg_file[94]), .ZN(n3177) );
  NAND4_X1 U3198 ( .A1(n6363), .A2(n6364), .A3(n3176), .A4(n3177), .ZN(n3178)
         );
  AOI22_X1 U3199 ( .A1(n3388), .A2(n3175), .B1(n6373), .B2(n3178), .ZN(n3179)
         );
  AOI22_X1 U3200 ( .A1(n3386), .A2(reg_file[414]), .B1(n3293), .B2(
        reg_file[510]), .ZN(n3180) );
  AOI22_X1 U3201 ( .A1(n4801), .A2(reg_file[478]), .B1(n4797), .B2(
        reg_file[446]), .ZN(n3181) );
  AOI22_X1 U3202 ( .A1(n4806), .A2(reg_file[350]), .B1(n3285), .B2(
        reg_file[382]), .ZN(n3182) );
  AOI22_X1 U3203 ( .A1(n4811), .A2(reg_file[286]), .B1(n4809), .B2(
        reg_file[318]), .ZN(n3183) );
  NAND4_X1 U3204 ( .A1(n3180), .A2(n3181), .A3(n3182), .A4(n3183), .ZN(n3184)
         );
  NAND4_X1 U3205 ( .A1(n6365), .A2(n6366), .A3(n6367), .A4(n6368), .ZN(n3185)
         );
  AOI22_X1 U3206 ( .A1(n3387), .A2(n3184), .B1(n3362), .B2(n3185), .ZN(n3186)
         );
  NAND2_X1 U3207 ( .A1(n3179), .A2(n3186), .ZN(rs1_val_gpr_w[30]) );
  OAI22_X1 U3208 ( .A1(reset_vector_i[5]), .A2(reset_vector_i[4]), .B1(
        n_0_net__4_), .B2(n6715), .ZN(n3187) );
  NOR2_X1 U3209 ( .A1(n3187), .A2(n6551), .ZN(n3188) );
  AOI21_X1 U3210 ( .B1(n3319), .B2(csr_mepc_w[5]), .A(n3188), .ZN(n3189) );
  AOI22_X1 U3211 ( .A1(reset_vector_i[5]), .A2(n6554), .B1(mem_i_pc_o[5]), 
        .B2(n6588), .ZN(n3190) );
  XOR2_X1 U3212 ( .A(DP_OP_181_135_5161_n28), .B(DP_OP_181_135_5161_n74), .Z(
        n3191) );
  NAND2_X1 U3213 ( .A1(DP_OP_181_135_5161_n95), .A2(n3191), .ZN(n3192) );
  OAI211_X1 U3214 ( .C1(DP_OP_181_135_5161_n95), .C2(n3191), .A(n6559), .B(
        n3192), .ZN(n3193) );
  NAND3_X1 U3215 ( .A1(n3189), .A2(n3190), .A3(n3193), .ZN(n2911) );
  AOI22_X1 U3216 ( .A1(n3355), .A2(reg_file[668]), .B1(n3293), .B2(
        reg_file[764]), .ZN(n3194) );
  AOI22_X1 U3217 ( .A1(n4796), .A2(reg_file[700]), .B1(n4800), .B2(
        reg_file[732]), .ZN(n3195) );
  AOI22_X1 U3218 ( .A1(n3286), .A2(reg_file[636]), .B1(n4805), .B2(
        reg_file[604]), .ZN(n3196) );
  AOI22_X1 U3219 ( .A1(n4807), .A2(reg_file[572]), .B1(n4812), .B2(
        reg_file[540]), .ZN(n3197) );
  NAND4_X1 U3220 ( .A1(n3194), .A2(n3195), .A3(n3196), .A4(n3197), .ZN(n3198)
         );
  AOI22_X1 U3221 ( .A1(n4813), .A2(reg_file[508]), .B1(n3386), .B2(
        reg_file[412]), .ZN(n3199) );
  AOI22_X1 U3222 ( .A1(n4796), .A2(reg_file[444]), .B1(n4801), .B2(
        reg_file[476]), .ZN(n3200) );
  AOI22_X1 U3223 ( .A1(n3285), .A2(reg_file[380]), .B1(n4806), .B2(
        reg_file[348]), .ZN(n3201) );
  AOI22_X1 U3224 ( .A1(n4809), .A2(reg_file[316]), .B1(n4811), .B2(
        reg_file[284]), .ZN(n3202) );
  NAND4_X1 U3225 ( .A1(n3199), .A2(n3200), .A3(n3201), .A4(n3202), .ZN(n3203)
         );
  AOI22_X1 U3226 ( .A1(n3388), .A2(n3198), .B1(n3387), .B2(n3203), .ZN(n3204)
         );
  AOI22_X1 U3227 ( .A1(n3293), .A2(reg_file[1020]), .B1(n4790), .B2(
        reg_file[924]), .ZN(n3205) );
  AOI22_X1 U3228 ( .A1(n4796), .A2(reg_file[956]), .B1(n4801), .B2(
        reg_file[988]), .ZN(n3206) );
  AOI22_X1 U3229 ( .A1(n3285), .A2(reg_file[892]), .B1(n4806), .B2(
        reg_file[860]), .ZN(n3207) );
  AOI22_X1 U3230 ( .A1(n4809), .A2(reg_file[828]), .B1(n4811), .B2(
        reg_file[796]), .ZN(n3208) );
  NAND4_X1 U3231 ( .A1(n3205), .A2(n3206), .A3(n3207), .A4(n3208), .ZN(n3209)
         );
  AOI22_X1 U3232 ( .A1(n3386), .A2(reg_file[156]), .B1(n4814), .B2(
        reg_file[252]), .ZN(n3210) );
  AOI22_X1 U3233 ( .A1(n4796), .A2(reg_file[188]), .B1(n4801), .B2(
        reg_file[220]), .ZN(n3211) );
  AOI22_X1 U3234 ( .A1(n3286), .A2(reg_file[124]), .B1(n4806), .B2(
        reg_file[92]), .ZN(n3212) );
  AOI22_X1 U3235 ( .A1(n4809), .A2(reg_file[60]), .B1(n4812), .B2(reg_file[28]), .ZN(n3213) );
  NAND4_X1 U3236 ( .A1(n3210), .A2(n3211), .A3(n3212), .A4(n3213), .ZN(n3214)
         );
  AOI22_X1 U3237 ( .A1(n3362), .A2(n3209), .B1(n6373), .B2(n3214), .ZN(n3215)
         );
  NAND2_X2 U3238 ( .A1(n3204), .A2(n3215), .ZN(rs1_val_gpr_w[28]) );
  INV_X1 U3239 ( .A(reset_vector_i[18]), .ZN(n3216) );
  INV_X1 U3240 ( .A(n6697), .ZN(n3217) );
  AOI221_X1 U3241 ( .B1(reset_vector_i[18]), .B2(n6697), .C1(n3216), .C2(n3217), .A(n6551), .ZN(n3218) );
  AOI21_X1 U3242 ( .B1(n3319), .B2(csr_mepc_w[18]), .A(n3218), .ZN(n3219) );
  AOI22_X1 U3243 ( .A1(reset_vector_i[18]), .A2(n6554), .B1(mem_i_pc_o[18]), 
        .B2(n6588), .ZN(n3220) );
  XNOR2_X1 U3244 ( .A(n3430), .B(DP_OP_181_135_5161_n108), .ZN(n3221) );
  NAND2_X1 U3245 ( .A1(DP_OP_181_135_5161_n87), .A2(n3221), .ZN(n3222) );
  OAI211_X1 U3246 ( .C1(DP_OP_181_135_5161_n87), .C2(n3221), .A(n3363), .B(
        n3222), .ZN(n3223) );
  NAND3_X1 U3247 ( .A1(n3219), .A2(n3220), .A3(n3223), .ZN(n2898) );
  INV_X1 U3248 ( .A(reset_vector_i[1]), .ZN(n3224) );
  AOI22_X1 U3249 ( .A1(mem_i_pc_o[1]), .A2(n6588), .B1(csr_mepc_w[1]), .B2(
        n3319), .ZN(n3225) );
  XOR2_X1 U3250 ( .A(DP_OP_181_135_5161_n70), .B(DP_OP_181_135_5161_n32), .Z(
        n3226) );
  NAND2_X1 U3251 ( .A1(DP_OP_181_135_5161_n91), .A2(n3226), .ZN(n3227) );
  OAI211_X1 U3252 ( .C1(DP_OP_181_135_5161_n91), .C2(n3226), .A(n3363), .B(
        n3227), .ZN(n3228) );
  OAI211_X1 U3253 ( .C1(n6593), .C2(n3224), .A(n3225), .B(n3228), .ZN(n2915)
         );
  INV_X1 U3254 ( .A(sub_x_59_n28), .ZN(n3229) );
  OAI21_X1 U3255 ( .B1(rs1_val_gpr_w[16]), .B2(n3338), .A(n3229), .ZN(n3513)
         );
  OAI21_X1 U3256 ( .B1(n3379), .B2(rs2_val_gpr_w[6]), .A(n3558), .ZN(n3530) );
  AND3_X1 U3257 ( .A1(n3556), .A2(rs2_val_gpr_w[10]), .A3(n3525), .ZN(n3230)
         );
  AOI21_X1 U3258 ( .B1(n3289), .B2(rs2_val_gpr_w[11]), .A(n3230), .ZN(n3537)
         );
  NOR2_X1 U3259 ( .A1(n3648), .A2(n3542), .ZN(n3231) );
  NOR3_X1 U3260 ( .A1(n3648), .A2(n3518), .A3(n3517), .ZN(n3232) );
  AOI211_X1 U3261 ( .C1(n3349), .C2(rs2_val_gpr_w[19]), .A(n3231), .B(n3232), 
        .ZN(n3516) );
  NAND2_X1 U3262 ( .A1(n3333), .A2(rs2_val_gpr_w[26]), .ZN(n3233) );
  NAND2_X1 U3263 ( .A1(n3331), .A2(rs2_val_gpr_w[27]), .ZN(n3234) );
  OAI21_X1 U3264 ( .B1(n3233), .B2(n3662), .A(n3234), .ZN(n3235) );
  AOI22_X1 U3265 ( .A1(n3320), .A2(rs2_val_gpr_w[28]), .B1(n3481), .B2(n3235), 
        .ZN(n3236) );
  NOR2_X1 U3266 ( .A1(n3236), .A2(n3460), .ZN(n3237) );
  AOI21_X1 U3267 ( .B1(rs2_val_gpr_w[29]), .B2(n3305), .A(n3237), .ZN(n3399)
         );
  AOI21_X1 U3268 ( .B1(sub_x_59_n1), .B2(n3406), .A(n3404), .ZN(n3238) );
  NAND2_X1 U3269 ( .A1(n3470), .A2(n3238), .ZN(n3401) );
  INV_X1 U3270 ( .A(n3424), .ZN(n3239) );
  NOR2_X1 U3271 ( .A1(n3423), .A2(n3239), .ZN(n3396) );
  INV_X1 U3272 ( .A(n6413), .ZN(n3240) );
  INV_X1 U3273 ( .A(n6853), .ZN(n3241) );
  OAI21_X1 U3274 ( .B1(n3240), .B2(n6854), .A(n6855), .ZN(n3242) );
  NAND2_X1 U3275 ( .A1(n3242), .A2(n3241), .ZN(n6866) );
  AOI22_X1 U3276 ( .A1(n4756), .A2(reg_file[729]), .B1(n4758), .B2(
        reg_file[761]), .ZN(n3243) );
  AOI22_X1 U3277 ( .A1(n4767), .A2(reg_file[665]), .B1(n4818), .B2(
        reg_file[697]), .ZN(n3244) );
  AOI22_X1 U3278 ( .A1(n3799), .A2(reg_file[601]), .B1(n4780), .B2(
        reg_file[633]), .ZN(n3245) );
  AOI22_X1 U3279 ( .A1(n4788), .A2(reg_file[537]), .B1(n4786), .B2(
        reg_file[569]), .ZN(n3246) );
  NAND4_X1 U3280 ( .A1(n3243), .A2(n3244), .A3(n3245), .A4(n3246), .ZN(n3247)
         );
  AOI22_X1 U3281 ( .A1(n4758), .A2(reg_file[505]), .B1(n3519), .B2(
        reg_file[473]), .ZN(n3248) );
  AOI22_X1 U3282 ( .A1(n4767), .A2(reg_file[409]), .B1(n4818), .B2(
        reg_file[441]), .ZN(n3249) );
  AOI22_X1 U3283 ( .A1(n3799), .A2(reg_file[345]), .B1(n4780), .B2(
        reg_file[377]), .ZN(n3250) );
  AOI22_X1 U3284 ( .A1(n4788), .A2(reg_file[281]), .B1(n4787), .B2(
        reg_file[313]), .ZN(n3251) );
  NAND4_X1 U3285 ( .A1(n3248), .A2(n3249), .A3(n3250), .A4(n3251), .ZN(n3252)
         );
  AOI22_X1 U3286 ( .A1(n5808), .A2(n3247), .B1(n5804), .B2(n3252), .ZN(n3253)
         );
  AOI22_X1 U3287 ( .A1(n4758), .A2(reg_file[249]), .B1(n4757), .B2(
        reg_file[217]), .ZN(n3254) );
  AOI22_X1 U3288 ( .A1(n4767), .A2(reg_file[153]), .B1(n4818), .B2(
        reg_file[185]), .ZN(n3255) );
  AOI22_X1 U3289 ( .A1(n3799), .A2(reg_file[89]), .B1(n4779), .B2(
        reg_file[121]), .ZN(n3256) );
  AOI22_X1 U3290 ( .A1(n4788), .A2(reg_file[25]), .B1(n4787), .B2(reg_file[57]), .ZN(n3257) );
  NAND4_X1 U3291 ( .A1(n3254), .A2(n3255), .A3(n3256), .A4(n3257), .ZN(n3258)
         );
  AOI22_X1 U3292 ( .A1(n4758), .A2(reg_file[1017]), .B1(n4755), .B2(
        reg_file[985]), .ZN(n3259) );
  AOI22_X1 U3293 ( .A1(n4767), .A2(reg_file[921]), .B1(n4818), .B2(
        reg_file[953]), .ZN(n3260) );
  AOI22_X1 U3294 ( .A1(n3799), .A2(reg_file[857]), .B1(n4779), .B2(
        reg_file[889]), .ZN(n3261) );
  AOI22_X1 U3295 ( .A1(n4788), .A2(reg_file[793]), .B1(n4787), .B2(
        reg_file[825]), .ZN(n3262) );
  NAND4_X1 U3296 ( .A1(n3259), .A2(n3260), .A3(n3261), .A4(n3262), .ZN(n3263)
         );
  AOI22_X1 U3297 ( .A1(n5805), .A2(n3258), .B1(n4816), .B2(n3263), .ZN(n3264)
         );
  NAND2_X1 U3298 ( .A1(n3253), .A2(n3264), .ZN(rs2_val_gpr_w[25]) );
  NAND4_X1 U3299 ( .A1(n5914), .A2(n5915), .A3(n5916), .A4(n5917), .ZN(n3265)
         );
  NAND4_X1 U3300 ( .A1(n5918), .A2(n5919), .A3(n5920), .A4(n5921), .ZN(n3266)
         );
  AOI22_X1 U3301 ( .A1(n6381), .A2(n3265), .B1(n3362), .B2(n3266), .ZN(n3267)
         );
  NAND4_X1 U3302 ( .A1(n5927), .A2(n5928), .A3(n5929), .A4(n5930), .ZN(n3268)
         );
  AOI22_X1 U3303 ( .A1(n6373), .A2(n5926), .B1(n6392), .B2(n3268), .ZN(n3269)
         );
  NAND2_X1 U3304 ( .A1(n3267), .A2(n3269), .ZN(rs1_val_gpr_w[5]) );
  INV_X1 U3305 ( .A(reset_vector_i[14]), .ZN(n3270) );
  INV_X1 U3306 ( .A(n6703), .ZN(n3271) );
  AOI221_X1 U3307 ( .B1(reset_vector_i[14]), .B2(n6703), .C1(n3270), .C2(n3271), .A(n6551), .ZN(n3272) );
  AOI21_X1 U3308 ( .B1(n3319), .B2(csr_mepc_w[14]), .A(n3272), .ZN(n3273) );
  AOI22_X1 U3309 ( .A1(reset_vector_i[14]), .A2(n6554), .B1(mem_i_pc_o[14]), 
        .B2(n6588), .ZN(n3274) );
  XNOR2_X1 U3310 ( .A(n3419), .B(DP_OP_181_135_5161_n104), .ZN(n3275) );
  NAND2_X1 U3311 ( .A1(DP_OP_181_135_5161_n83), .A2(n3275), .ZN(n3276) );
  OAI211_X1 U3312 ( .C1(DP_OP_181_135_5161_n83), .C2(n3275), .A(n3363), .B(
        n3276), .ZN(n3277) );
  NAND3_X1 U3313 ( .A1(n3273), .A2(n3274), .A3(n3277), .ZN(n2902) );
  INV_X1 U3314 ( .A(reset_vector_i[2]), .ZN(n3278) );
  AOI22_X1 U3315 ( .A1(mem_i_pc_o[2]), .A2(n6588), .B1(csr_mepc_w[2]), .B2(
        n3319), .ZN(n3279) );
  XNOR2_X1 U3316 ( .A(n3450), .B(DP_OP_181_135_5161_n92), .ZN(n3280) );
  NAND2_X1 U3317 ( .A1(C1_Z_2), .A2(n3280), .ZN(n3281) );
  OAI211_X1 U3318 ( .C1(C1_Z_2), .C2(n3280), .A(n3363), .B(n3281), .ZN(n3282)
         );
  OAI211_X1 U3319 ( .C1(n6593), .C2(n3278), .A(n3279), .B(n3282), .ZN(n2914)
         );
  NAND2_X1 U3320 ( .A1(n6788), .A2(n6789), .ZN(n3283) );
  AOI221_X1 U3321 ( .B1(muldiv_ready_w), .B2(rd_wr_en_q), .C1(n6786), .C2(
        rd_wr_en_q), .A(rst_i), .ZN(n3284) );
  OAI22_X1 U3322 ( .A1(n6787), .A2(n3283), .B1(n6813), .B2(n3284), .ZN(n2875)
         );
  BUF_X4 U3323 ( .A(n5813), .Z(n4788) );
  BUF_X4 U3324 ( .A(n5810), .Z(n4758) );
  BUF_X2 U3325 ( .A(n5810), .Z(n4759) );
  BUF_X2 U3326 ( .A(n6387), .Z(n4812) );
  BUF_X2 U3327 ( .A(n6387), .Z(n4811) );
  INV_X4 U3328 ( .A(n6586), .ZN(n3297) );
  BUF_X4 U3329 ( .A(n6386), .Z(n4809) );
  BUF_X2 U3330 ( .A(n6386), .Z(n4807) );
  BUF_X2 U3331 ( .A(n6386), .Z(n4808) );
  BUF_X2 U3332 ( .A(n6384), .Z(n4800) );
  BUF_X2 U3333 ( .A(n6384), .Z(n4798) );
  BUF_X2 U3334 ( .A(n6384), .Z(n4801) );
  BUF_X4 U3335 ( .A(n5812), .Z(n4787) );
  BUF_X2 U3336 ( .A(n5812), .Z(n4786) );
  AND2_X2 U3337 ( .A1(n6400), .A2(mem_i_inst_i[20]), .ZN(n5809) );
  BUF_X2 U3338 ( .A(n5809), .Z(n4756) );
  BUF_X4 U3339 ( .A(n5809), .Z(n4757) );
  BUF_X2 U3340 ( .A(n6382), .Z(n3386) );
  BUF_X4 U3341 ( .A(n6382), .Z(n3355) );
  NOR2_X1 U3342 ( .A1(n4942), .A2(n6608), .ZN(n6382) );
  AND2_X2 U3343 ( .A1(n4943), .A2(n6608), .ZN(n6396) );
  BUF_X4 U3344 ( .A(n6396), .Z(n4815) );
  INV_X2 U3345 ( .A(n4820), .ZN(n4819) );
  OR2_X2 U3346 ( .A1(n6466), .A2(n6579), .ZN(n4820) );
  NAND4_X2 U3347 ( .A1(n5841), .A2(n5840), .A3(n5839), .A4(n5838), .ZN(
        rs1_val_gpr_w[1]) );
  BUF_X8 U3348 ( .A(n3768), .Z(n3285) );
  BUF_X8 U3349 ( .A(n3768), .Z(n3286) );
  NAND4_X2 U3350 ( .A1(n5865), .A2(n5862), .A3(n5863), .A4(n5864), .ZN(
        rs1_val_gpr_w[2]) );
  INV_X1 U3351 ( .A(n4820), .ZN(n3287) );
  NAND2_X1 U3352 ( .A1(rs2_val_gpr_w[18]), .A2(n3334), .ZN(n3542) );
  NAND2_X1 U3353 ( .A1(n3338), .A2(rs1_val_gpr_w[16]), .ZN(n3578) );
  NAND4_X1 U3354 ( .A1(n6098), .A2(n6097), .A3(n6096), .A4(n6095), .ZN(
        rs1_val_gpr_w[12]) );
  INV_X1 U3355 ( .A(rs1_val_gpr_w[3]), .ZN(n3288) );
  NAND4_X2 U3356 ( .A1(n5057), .A2(n5056), .A3(n5055), .A4(n5054), .ZN(
        rs2_val_gpr_w[1]) );
  NAND4_X1 U3357 ( .A1(n5114), .A2(n5113), .A3(n5112), .A4(n5111), .ZN(
        rs2_val_gpr_w[2]) );
  NAND4_X1 U3358 ( .A1(n5170), .A2(n5169), .A3(n5168), .A4(n5167), .ZN(
        rs2_val_gpr_w[3]) );
  NAND4_X1 U3359 ( .A1(n6002), .A2(n6001), .A3(n6000), .A4(n5999), .ZN(
        rs1_val_gpr_w[8]) );
  INV_X1 U3360 ( .A(rs1_val_gpr_w[11]), .ZN(n3289) );
  NAND4_X1 U3361 ( .A1(n6026), .A2(n6025), .A3(n6024), .A4(n6023), .ZN(
        rs1_val_gpr_w[9]) );
  INV_X1 U3362 ( .A(rs1_val_gpr_w[13]), .ZN(n3290) );
  NAND4_X1 U3363 ( .A1(n6204), .A2(n6203), .A3(n6202), .A4(n6201), .ZN(
        rs1_val_gpr_w[17]) );
  NAND4_X1 U3364 ( .A1(n6228), .A2(n6227), .A3(n6226), .A4(n6225), .ZN(
        rs1_val_gpr_w[18]) );
  NAND4_X1 U3365 ( .A1(n5913), .A2(n5912), .A3(n5911), .A4(n5910), .ZN(
        rs1_val_gpr_w[4]) );
  NAND4_X1 U3366 ( .A1(n5659), .A2(n5658), .A3(n5657), .A4(n5656), .ZN(
        rs2_val_gpr_w[23]) );
  INV_X1 U3367 ( .A(rs2_val_gpr_w[13]), .ZN(n3291) );
  INV_X1 U3368 ( .A(rs2_val_gpr_w[7]), .ZN(n3292) );
  INV_X1 U3369 ( .A(n6918), .ZN(n4827) );
  INV_X1 U3370 ( .A(n7867), .ZN(n7802) );
  INV_X1 U3371 ( .A(n3317), .ZN(n4814) );
  BUF_X1 U3372 ( .A(n6384), .Z(n3314) );
  BUF_X1 U3373 ( .A(n6387), .Z(n3316) );
  BUF_X1 U3374 ( .A(n6386), .Z(n3315) );
  BUF_X1 U3375 ( .A(n5812), .Z(n3318) );
  INV_X2 U3376 ( .A(n3317), .ZN(n3293) );
  BUF_X4 U3377 ( .A(n6404), .Z(n3294) );
  AND2_X1 U3378 ( .A1(n4943), .A2(mem_i_inst_i[16]), .ZN(n6383) );
  BUF_X2 U3379 ( .A(n6385), .Z(n3295) );
  BUF_X2 U3380 ( .A(n5813), .Z(n3296) );
  AND2_X2 U3381 ( .A1(n6400), .A2(n6623), .ZN(n5810) );
  AND3_X2 U3382 ( .A1(n6410), .A2(mem_i_inst_i[21]), .A3(mem_i_inst_i[20]), 
        .ZN(n3769) );
  AND2_X2 U3383 ( .A1(n4975), .A2(mem_i_inst_i[22]), .ZN(n5811) );
  AND3_X2 U3384 ( .A1(n6411), .A2(mem_i_inst_i[20]), .A3(mem_i_inst_i[22]), 
        .ZN(n3799) );
  AND2_X1 U3385 ( .A1(mem_i_inst_i[24]), .A2(mem_i_inst_i[23]), .ZN(n5805) );
  AND2_X2 U3386 ( .A1(mem_i_inst_i[19]), .A2(mem_i_inst_i[18]), .ZN(n6373) );
  BUF_X1 U3387 ( .A(n6559), .Z(n3363) );
  NAND2_X1 U3388 ( .A1(n6465), .A2(n6463), .ZN(n6581) );
  INV_X1 U3389 ( .A(n6551), .ZN(n6555) );
  NOR2_X1 U3390 ( .A1(rs2_val_gpr_w[14]), .A2(n3323), .ZN(n3554) );
  NAND2_X1 U3391 ( .A1(rs2_val_gpr_w[8]), .A2(n3321), .ZN(n3544) );
  NAND2_X1 U3392 ( .A1(rs2_val_gpr_w[20]), .A2(n3341), .ZN(n3540) );
  NOR2_X1 U3393 ( .A1(rs2_val_gpr_w[20]), .A2(n3341), .ZN(n3549) );
  NAND2_X1 U3394 ( .A1(n3350), .A2(rs1_val_gpr_w[12]), .ZN(n3584) );
  NOR2_X1 U3395 ( .A1(n3343), .A2(rs1_val_gpr_w[22]), .ZN(n3510) );
  NAND2_X1 U3396 ( .A1(n3378), .A2(rs1_val_gpr_w[14]), .ZN(n3581) );
  NAND2_X1 U3397 ( .A1(n3382), .A2(rs1_val_gpr_w[8]), .ZN(n3582) );
  INV_X1 U3398 ( .A(n3526), .ZN(n3521) );
  AND2_X1 U3399 ( .A1(n3343), .A2(rs1_val_gpr_w[22]), .ZN(n3509) );
  INV_X1 U3400 ( .A(rs2_val_gpr_w[31]), .ZN(n3298) );
  INV_X1 U3401 ( .A(rs2_val_gpr_w[3]), .ZN(n3299) );
  INV_X1 U3402 ( .A(rs1_val_gpr_w[17]), .ZN(n3300) );
  NAND4_X2 U3403 ( .A1(n6122), .A2(n6121), .A3(n6120), .A4(n6119), .ZN(
        rs1_val_gpr_w[13]) );
  INV_X1 U3404 ( .A(rs1_val_gpr_w[21]), .ZN(n3301) );
  NAND4_X1 U3405 ( .A1(n5889), .A2(n5888), .A3(n5887), .A4(n5886), .ZN(
        rs1_val_gpr_w[3]) );
  INV_X1 U3406 ( .A(rs2_val_gpr_w[1]), .ZN(n3302) );
  NAND4_X1 U3407 ( .A1(n5000), .A2(n4999), .A3(n4998), .A4(n4997), .ZN(
        rs2_val_gpr_w[0]) );
  INV_X1 U3408 ( .A(rs2_val_gpr_w[5]), .ZN(n3303) );
  INV_X1 U3409 ( .A(rs1_val_gpr_w[15]), .ZN(n3304) );
  NAND4_X2 U3410 ( .A1(n6074), .A2(n6072), .A3(n6073), .A4(n6071), .ZN(
        rs1_val_gpr_w[11]) );
  INV_X1 U3411 ( .A(rs1_val_gpr_w[29]), .ZN(n3305) );
  INV_X1 U3412 ( .A(rs1_val_gpr_w[5]), .ZN(n3306) );
  INV_X1 U3413 ( .A(rs1_val_gpr_w[23]), .ZN(n3307) );
  INV_X1 U3414 ( .A(rs1_val_gpr_w[9]), .ZN(n3308) );
  NAND4_X1 U3415 ( .A1(n5954), .A2(n5953), .A3(n5952), .A4(n5951), .ZN(
        rs1_val_gpr_w[6]) );
  NAND4_X1 U3416 ( .A1(n5978), .A2(n5977), .A3(n5976), .A4(n5975), .ZN(
        rs1_val_gpr_w[7]) );
  INV_X1 U3417 ( .A(rs2_val_gpr_w[2]), .ZN(n3309) );
  INV_X1 U3418 ( .A(rs2_val_gpr_w[23]), .ZN(n3310) );
  INV_X1 U3419 ( .A(rs2_val_gpr_w[15]), .ZN(n3311) );
  NAND4_X1 U3420 ( .A1(n5363), .A2(n5362), .A3(n5361), .A4(n5360), .ZN(
        rs2_val_gpr_w[9]) );
  INV_X1 U3421 ( .A(rs2_val_gpr_w[21]), .ZN(n3312) );
  NAND4_X1 U3422 ( .A1(n5339), .A2(n5338), .A3(n5337), .A4(n5336), .ZN(
        rs2_val_gpr_w[8]) );
  NAND4_X1 U3423 ( .A1(n5315), .A2(n5314), .A3(n5313), .A4(n5312), .ZN(
        rs2_val_gpr_w[7]) );
  NAND4_X1 U3424 ( .A1(n5406), .A2(n5405), .A3(n5404), .A4(n5403), .ZN(
        rs2_val_gpr_w[11]) );
  INV_X1 U3425 ( .A(rs2_val_gpr_w[6]), .ZN(n3313) );
  INV_X1 U3426 ( .A(n4817), .ZN(n3357) );
  BUF_X1 U3427 ( .A(n6384), .Z(n3356) );
  BUF_X1 U3428 ( .A(n6387), .Z(n3358) );
  BUF_X1 U3429 ( .A(n6383), .Z(n3360) );
  NOR2_X1 U3430 ( .A1(n6619), .A2(mem_i_inst_i[18]), .ZN(n6381) );
  INV_X1 U3431 ( .A(n3800), .ZN(n3361) );
  INV_X1 U3432 ( .A(n6396), .ZN(n3317) );
  NOR2_X1 U3433 ( .A1(n6615), .A2(mem_i_inst_i[19]), .ZN(n6392) );
  AND3_X2 U3434 ( .A1(n6608), .A2(n6604), .A3(mem_i_inst_i[17]), .ZN(n3768) );
  NAND2_X1 U3435 ( .A1(mem_i_inst_i[16]), .A2(mem_i_inst_i[17]), .ZN(n4945) );
  NOR2_X1 U3436 ( .A1(mem_i_inst_i[21]), .A2(mem_i_inst_i[22]), .ZN(n6400) );
  OAI21_X1 U3437 ( .B1(n3423), .B2(n3395), .A(n3422), .ZN(n3394) );
  NAND2_X1 U3438 ( .A1(n3486), .A2(n3435), .ZN(n3485) );
  NOR3_X1 U3439 ( .A1(n7826), .A2(n7825), .A3(n7824), .ZN(n7827) );
  XNOR2_X1 U3440 ( .A(DP_OP_181_135_5161_n117), .B(n3435), .ZN(n3443) );
  BUF_X2 U3441 ( .A(n7794), .Z(n3364) );
  NOR3_X1 U3442 ( .A1(n7695), .A2(n7694), .A3(n7693), .ZN(n7696) );
  AND4_X2 U3443 ( .A1(n7727), .A2(n7726), .A3(n7725), .A4(n7724), .ZN(n7728)
         );
  BUF_X2 U3444 ( .A(n7614), .Z(n3365) );
  BUF_X2 U3445 ( .A(n7567), .Z(n3366) );
  AND2_X1 U3446 ( .A1(n3425), .A2(n3416), .ZN(n3415) );
  INV_X1 U3447 ( .A(n6577), .ZN(n6583) );
  BUF_X2 U3448 ( .A(n6589), .Z(n3319) );
  BUF_X1 U3449 ( .A(n7137), .Z(n3371) );
  XNOR2_X1 U3450 ( .A(rs1_val_gpr_w[31]), .B(rs2_val_gpr_w[31]), .ZN(
        sub_x_60_n1) );
  OR2_X1 U3451 ( .A1(n3384), .A2(rs1_val_gpr_w[25]), .ZN(n3499) );
  NAND2_X1 U3452 ( .A1(n3384), .A2(rs1_val_gpr_w[25]), .ZN(n3497) );
  OR2_X1 U3453 ( .A1(n3385), .A2(rs1_val_gpr_w[26]), .ZN(n3487) );
  OR2_X1 U3454 ( .A1(n3376), .A2(rs1_val_gpr_w[27]), .ZN(n3488) );
  INV_X1 U3455 ( .A(n3525), .ZN(rs1_val_gpr_w[10]) );
  INV_X1 U3456 ( .A(rs1_val_gpr_w[28]), .ZN(n3320) );
  INV_X1 U3457 ( .A(rs1_val_gpr_w[8]), .ZN(n3321) );
  INV_X1 U3458 ( .A(rs2_val_gpr_w[11]), .ZN(n3322) );
  INV_X1 U3459 ( .A(rs1_val_gpr_w[14]), .ZN(n3323) );
  INV_X1 U3460 ( .A(rs1_val_gpr_w[4]), .ZN(n3324) );
  INV_X1 U3461 ( .A(rs2_val_gpr_w[4]), .ZN(n3325) );
  INV_X1 U3462 ( .A(rs2_val_gpr_w[20]), .ZN(n3326) );
  INV_X1 U3463 ( .A(rs1_val_gpr_w[7]), .ZN(n3327) );
  INV_X1 U3464 ( .A(rs2_val_gpr_w[0]), .ZN(n3328) );
  INV_X1 U3465 ( .A(rs1_val_gpr_w[2]), .ZN(n3329) );
  INV_X1 U3466 ( .A(rs1_val_gpr_w[25]), .ZN(n3330) );
  INV_X1 U3467 ( .A(rs1_val_gpr_w[27]), .ZN(n3331) );
  INV_X1 U3468 ( .A(rs2_val_gpr_w[19]), .ZN(n3332) );
  INV_X1 U3469 ( .A(rs1_val_gpr_w[26]), .ZN(n3333) );
  INV_X1 U3470 ( .A(rs1_val_gpr_w[18]), .ZN(n3334) );
  INV_X1 U3471 ( .A(rs1_val_gpr_w[24]), .ZN(n3335) );
  INV_X1 U3472 ( .A(rs2_val_gpr_w[24]), .ZN(n3336) );
  INV_X1 U3473 ( .A(rs2_val_gpr_w[18]), .ZN(n3337) );
  INV_X1 U3474 ( .A(rs2_val_gpr_w[16]), .ZN(n3338) );
  INV_X1 U3475 ( .A(rs1_val_gpr_w[16]), .ZN(n3339) );
  INV_X1 U3476 ( .A(rs2_val_gpr_w[17]), .ZN(n3340) );
  INV_X1 U3477 ( .A(rs1_val_gpr_w[20]), .ZN(n3341) );
  INV_X1 U3478 ( .A(rs2_val_gpr_w[29]), .ZN(n3342) );
  INV_X1 U3479 ( .A(rs2_val_gpr_w[22]), .ZN(n3343) );
  INV_X1 U3480 ( .A(rs1_val_gpr_w[22]), .ZN(n3344) );
  INV_X1 U3481 ( .A(rs1_val_gpr_w[31]), .ZN(n3345) );
  INV_X1 U3482 ( .A(rs2_val_gpr_w[30]), .ZN(n3346) );
  INV_X1 U3483 ( .A(rs1_val_gpr_w[30]), .ZN(n3347) );
  INV_X1 U3484 ( .A(rs2_val_gpr_w[28]), .ZN(n3348) );
  INV_X1 U3485 ( .A(rs1_val_gpr_w[19]), .ZN(n3349) );
  INV_X1 U3486 ( .A(rs2_val_gpr_w[12]), .ZN(n3350) );
  INV_X1 U3487 ( .A(rs1_val_gpr_w[12]), .ZN(n3351) );
  BUF_X1 U3488 ( .A(n6382), .Z(n4790) );
  BUF_X1 U3489 ( .A(n6384), .Z(n4799) );
  INV_X2 U3490 ( .A(n3764), .ZN(n3352) );
  INV_X2 U3491 ( .A(n3842), .ZN(n3353) );
  BUF_X1 U3492 ( .A(n6385), .Z(n4806) );
  BUF_X1 U3493 ( .A(n5811), .Z(n4783) );
  BUF_X1 U3494 ( .A(n5813), .Z(n4789) );
  BUF_X2 U3495 ( .A(n6404), .Z(n4818) );
  BUF_X1 U3496 ( .A(n5808), .Z(n3390) );
  BUF_X1 U3497 ( .A(n5809), .Z(n4755) );
  BUF_X1 U3498 ( .A(n5804), .Z(n3389) );
  INV_X1 U3499 ( .A(n3317), .ZN(n3354) );
  BUF_X1 U3500 ( .A(n6392), .Z(n3388) );
  BUF_X1 U3501 ( .A(n6387), .Z(n4810) );
  BUF_X1 U3502 ( .A(n6381), .Z(n3387) );
  NOR2_X1 U3503 ( .A1(n4976), .A2(mem_i_inst_i[20]), .ZN(n5812) );
  AND2_X1 U3504 ( .A1(n4974), .A2(mem_i_inst_i[21]), .ZN(n6404) );
  BUF_X2 U3505 ( .A(n6385), .Z(n3359) );
  BUF_X2 U3506 ( .A(n6397), .Z(n3362) );
  XNOR2_X1 U3507 ( .A(DP_OP_181_135_5161_n3), .B(n3482), .ZN(
        U4_RSOP_173_C3_DATA1_30) );
  AOI21_X1 U3508 ( .B1(DP_OP_181_135_5161_n3), .B2(n3485), .A(n3484), .ZN(
        n3483) );
  XNOR2_X1 U3509 ( .A(n3444), .B(n3443), .ZN(U4_RSOP_173_C3_DATA1_27) );
  OAI21_X1 U3510 ( .B1(n3444), .B2(n3442), .A(n3441), .ZN(
        DP_OP_181_135_5161_n5) );
  AOI21_X1 U3511 ( .B1(DP_OP_181_135_5161_n7), .B2(n3446), .A(n3445), .ZN(
        n3444) );
  XNOR2_X1 U3512 ( .A(DP_OP_181_135_5161_n8), .B(n3440), .ZN(
        U4_RSOP_173_C3_DATA1_25) );
  XNOR2_X1 U3513 ( .A(DP_OP_181_135_5161_n7), .B(n3447), .ZN(
        U4_RSOP_173_C3_DATA1_26) );
  OAI22_X1 U3514 ( .A1(n3436), .A2(n3439), .B1(n3435), .B2(n3434), .ZN(
        DP_OP_181_135_5161_n7) );
  XNOR2_X1 U3515 ( .A(DP_OP_181_135_5161_n9), .B(n3438), .ZN(
        U4_RSOP_173_C3_DATA1_24) );
  OAI21_X1 U3516 ( .B1(n3430), .B2(n3429), .A(n3428), .ZN(
        DP_OP_181_135_5161_n14) );
  XNOR2_X1 U3517 ( .A(DP_OP_181_135_5161_n16), .B(n3433), .ZN(
        U4_RSOP_173_C3_DATA1_17) );
  AOI21_X1 U3518 ( .B1(DP_OP_181_135_5161_n16), .B2(n3432), .A(n3431), .ZN(
        n3430) );
  OAI21_X1 U3519 ( .B1(n3419), .B2(n3418), .A(n3417), .ZN(
        DP_OP_181_135_5161_n18) );
  XNOR2_X1 U3520 ( .A(DP_OP_181_135_5161_n20), .B(n3421), .ZN(
        U4_RSOP_173_C3_DATA1_13) );
  AOI22_X1 U3521 ( .A1(DP_OP_181_135_5161_n20), .A2(n3420), .B1(
        DP_OP_181_135_5161_n103), .B2(DP_OP_181_135_5161_n82), .ZN(n3419) );
  OAI21_X1 U3522 ( .B1(n3457), .B2(n3456), .A(n3455), .ZN(
        DP_OP_181_135_5161_n26) );
  AOI21_X1 U3523 ( .B1(DP_OP_181_135_5161_n28), .B2(n3459), .A(n3458), .ZN(
        n3457) );
  XNOR2_X1 U3524 ( .A(DP_OP_181_135_5161_n30), .B(n3496), .ZN(
        U4_RSOP_173_C3_DATA1_3) );
  BUF_X1 U3525 ( .A(n4973), .Z(n4753) );
  INV_X1 U3526 ( .A(n3394), .ZN(n3393) );
  BUF_X1 U3527 ( .A(n7827), .Z(n4844) );
  AOI21_X2 U3528 ( .B1(alu_a_q[0]), .B2(n7953), .A(n7952), .ZN(n4973) );
  OR2_X1 U3529 ( .A1(DP_OP_181_135_5161_n103), .A2(DP_OP_181_135_5161_n82), 
        .ZN(n3420) );
  INV_X1 U3530 ( .A(DP_OP_181_135_5161_n120), .ZN(n3486) );
  NOR2_X1 U3531 ( .A1(DP_OP_181_135_5161_n96), .A2(DP_OP_181_135_5161_n75), 
        .ZN(n3456) );
  NAND2_X1 U3532 ( .A1(DP_OP_181_135_5161_n96), .A2(DP_OP_181_135_5161_n75), 
        .ZN(n3455) );
  OR2_X1 U3533 ( .A1(DP_OP_181_135_5161_n95), .A2(DP_OP_181_135_5161_n74), 
        .ZN(n3459) );
  XNOR2_X1 U3534 ( .A(DP_OP_181_135_5161_n107), .B(DP_OP_181_135_5161_n86), 
        .ZN(n3433) );
  OR2_X1 U3535 ( .A1(DP_OP_181_135_5161_n107), .A2(DP_OP_181_135_5161_n86), 
        .ZN(n3432) );
  NAND2_X1 U3536 ( .A1(DP_OP_181_135_5161_n104), .A2(DP_OP_181_135_5161_n83), 
        .ZN(n3417) );
  NOR2_X1 U3537 ( .A1(DP_OP_181_135_5161_n100), .A2(DP_OP_181_135_5161_n79), 
        .ZN(n3423) );
  XNOR2_X1 U3538 ( .A(DP_OP_181_135_5161_n93), .B(DP_OP_181_135_5161_n72), 
        .ZN(n3496) );
  NOR2_X1 U3539 ( .A1(DP_OP_181_135_5161_n104), .A2(DP_OP_181_135_5161_n83), 
        .ZN(n3418) );
  NAND2_X1 U3540 ( .A1(DP_OP_181_135_5161_n99), .A2(DP_OP_181_135_5161_n78), 
        .ZN(n3395) );
  OR2_X1 U3541 ( .A1(DP_OP_181_135_5161_n99), .A2(DP_OP_181_135_5161_n78), 
        .ZN(n3424) );
  OR2_X1 U3542 ( .A1(DP_OP_181_135_5161_n116), .A2(n3391), .ZN(n3446) );
  NAND2_X1 U3543 ( .A1(DP_OP_181_135_5161_n93), .A2(DP_OP_181_135_5161_n72), 
        .ZN(n3492) );
  XNOR2_X1 U3544 ( .A(DP_OP_181_135_5161_n103), .B(DP_OP_181_135_5161_n82), 
        .ZN(n3421) );
  NAND2_X1 U3545 ( .A1(DP_OP_181_135_5161_n100), .A2(DP_OP_181_135_5161_n79), 
        .ZN(n3422) );
  NOR2_X1 U3546 ( .A1(DP_OP_181_135_5161_n108), .A2(DP_OP_181_135_5161_n87), 
        .ZN(n3429) );
  OR2_X1 U3547 ( .A1(DP_OP_181_135_5161_n114), .A2(DP_OP_181_135_5161_n89), 
        .ZN(n3437) );
  NAND2_X1 U3548 ( .A1(DP_OP_181_135_5161_n108), .A2(DP_OP_181_135_5161_n87), 
        .ZN(n3428) );
  BUF_X1 U3549 ( .A(n7863), .Z(n4845) );
  BUF_X1 U3550 ( .A(n7764), .Z(n4843) );
  OR2_X1 U3551 ( .A1(DP_OP_181_135_5161_n91), .A2(DP_OP_181_135_5161_n70), 
        .ZN(n3452) );
  AND2_X1 U3552 ( .A1(DP_OP_181_135_5161_n91), .A2(DP_OP_181_135_5161_n70), 
        .ZN(n3451) );
  AOI211_X1 U3553 ( .C1(n3352), .C2(n7862), .A(n7861), .B(n7860), .ZN(n7863)
         );
  BUF_X1 U3554 ( .A(n7696), .Z(n4842) );
  BUF_X1 U3555 ( .A(n7671), .Z(n4841) );
  AOI21_X1 U3556 ( .B1(n6579), .B2(mem_i_inst_i[31]), .A(n6561), .ZN(n6560) );
  OAI21_X1 U3557 ( .B1(n4718), .B2(n4715), .A(n4712), .ZN(n6579) );
  BUF_X1 U3558 ( .A(n7589), .Z(n4839) );
  BUF_X1 U3559 ( .A(n7545), .Z(n4838) );
  AOI21_X1 U3560 ( .B1(n7926), .B2(n7645), .A(n7927), .ZN(n7685) );
  BUF_X1 U3561 ( .A(n7520), .Z(n4837) );
  AOI22_X1 U3562 ( .A1(alu_a_q[22]), .A2(n3845), .B1(n7918), .B2(n7590), .ZN(
        n7628) );
  OR2_X1 U3563 ( .A1(n7921), .A2(n7576), .ZN(n7590) );
  INV_X1 U3564 ( .A(n7534), .ZN(n7555) );
  BUF_X2 U3565 ( .A(n7494), .Z(n3367) );
  OR2_X1 U3566 ( .A1(n6770), .A2(n6551), .ZN(n3453) );
  OAI21_X1 U3567 ( .B1(n7531), .B2(n7917), .A(n7914), .ZN(n7534) );
  BUF_X2 U3568 ( .A(n7404), .Z(n3368) );
  BUF_X2 U3569 ( .A(n7471), .Z(n3369) );
  AOI21_X1 U3570 ( .B1(alu_a_q[18]), .B2(n3838), .A(n7509), .ZN(n7531) );
  BUF_X1 U3571 ( .A(n7332), .Z(n4834) );
  BUF_X1 U3572 ( .A(n7365), .Z(n4835) );
  AND2_X1 U3573 ( .A1(n3501), .A2(n3500), .ZN(n3468) );
  BUF_X1 U3574 ( .A(n7275), .Z(n4832) );
  BUF_X1 U3575 ( .A(n7301), .Z(n4833) );
  OAI21_X1 U3576 ( .B1(n7890), .B2(n7458), .A(n7907), .ZN(n7460) );
  AOI22_X1 U3577 ( .A1(alu_a_q[18]), .A2(alu_b_q[18]), .B1(n7496), .B2(n7495), 
        .ZN(n7532) );
  OAI21_X1 U3578 ( .B1(n7408), .B2(n7905), .A(n7904), .ZN(n7458) );
  AOI22_X1 U3579 ( .A1(n3794), .A2(n3847), .B1(n7473), .B2(n7472), .ZN(n7496)
         );
  NOR2_X1 U3580 ( .A1(n7901), .A2(n7366), .ZN(n7408) );
  OAI21_X1 U3581 ( .B1(n3559), .B2(n3515), .A(n3511), .ZN(n3502) );
  OAI22_X1 U3582 ( .A1(alu_a_q[16]), .A2(alu_b_q[16]), .B1(n7444), .B2(n7443), 
        .ZN(n7472) );
  OAI22_X1 U3583 ( .A1(alu_a_q[13]), .A2(n3776), .B1(n7335), .B2(n7895), .ZN(
        n7366) );
  NOR2_X1 U3584 ( .A1(n7903), .A2(n7302), .ZN(n7335) );
  AOI22_X1 U3585 ( .A1(n3785), .A2(n3851), .B1(n7406), .B2(n7405), .ZN(n7443)
         );
  OAI22_X1 U3586 ( .A1(alu_a_q[14]), .A2(alu_b_q[14]), .B1(n7369), .B2(n7368), 
        .ZN(n7405) );
  OAI22_X1 U3587 ( .A1(alu_a_q[11]), .A2(n3775), .B1(n7291), .B2(n7897), .ZN(
        n7302) );
  BUF_X1 U3588 ( .A(n6845), .Z(n4821) );
  OAI21_X1 U3589 ( .B1(n3399), .B2(n3465), .A(n3464), .ZN(n3397) );
  AOI221_X1 U3590 ( .B1(n3776), .B2(n7337), .C1(n3815), .C2(n7337), .A(n7336), 
        .ZN(n7368) );
  OAI22_X1 U3591 ( .A1(alu_a_q[12]), .A2(alu_b_q[12]), .B1(n7304), .B2(n7303), 
        .ZN(n7337) );
  BUF_X2 U3592 ( .A(n7207), .Z(n3370) );
  OR2_X1 U3593 ( .A1(n3516), .A2(n3549), .ZN(n3508) );
  AND2_X1 U3594 ( .A1(n3408), .A2(n3409), .ZN(n3407) );
  AOI22_X1 U3595 ( .A1(n3408), .A2(n3405), .B1(sub_x_59_n1), .B2(n3409), .ZN(
        n3404) );
  AOI22_X1 U3596 ( .A1(n7240), .A2(n7239), .B1(n3811), .B2(alu_b_q[9]), .ZN(
        n7899) );
  INV_X1 U3597 ( .A(sub_x_59_n1), .ZN(n3408) );
  INV_X1 U3598 ( .A(n3410), .ZN(n3406) );
  NAND2_X1 U3599 ( .A1(n3410), .A2(n3409), .ZN(n3405) );
  AND3_X1 U3600 ( .A1(n3477), .A2(n3488), .A3(n3487), .ZN(n3414) );
  OAI22_X1 U3601 ( .A1(n7242), .A2(n7241), .B1(n3811), .B2(n3782), .ZN(n7252)
         );
  BUF_X2 U3602 ( .A(n7115), .Z(n3372) );
  INV_X1 U3603 ( .A(mem_addr_w[1]), .ZN(n6676) );
  AOI21_X1 U3604 ( .B1(sub_x_60_n28), .B2(n3541), .A(sub_x_60_n29), .ZN(n3518)
         );
  NOR2_X1 U3605 ( .A1(n3460), .A2(n3465), .ZN(n3398) );
  AOI22_X1 U3606 ( .A1(alu_a_q[8]), .A2(alu_b_q[8]), .B1(n7209), .B2(n7208), 
        .ZN(n7241) );
  BUF_X2 U3607 ( .A(n7093), .Z(n3373) );
  INV_X1 U3608 ( .A(n6740), .ZN(n3403) );
  INV_X1 U3609 ( .A(n3550), .ZN(n3517) );
  INV_X1 U3610 ( .A(mem_addr_w[0]), .ZN(n6673) );
  OR2_X1 U3611 ( .A1(n3320), .A2(rs2_val_gpr_w[28]), .ZN(n3481) );
  BUF_X2 U3612 ( .A(n5090), .Z(n3374) );
  OAI21_X1 U3613 ( .B1(n7188), .B2(n7187), .A(n7186), .ZN(n7208) );
  OR2_X1 U3614 ( .A1(n3342), .A2(rs1_val_gpr_w[29]), .ZN(n3471) );
  NOR2_X1 U3615 ( .A1(n3346), .A2(rs1_val_gpr_w[30]), .ZN(n3462) );
  NAND2_X1 U3616 ( .A1(n3310), .A2(rs1_val_gpr_w[23]), .ZN(n3500) );
  OR2_X1 U3617 ( .A1(n3348), .A2(rs1_val_gpr_w[28]), .ZN(n3477) );
  OR2_X1 U3618 ( .A1(n3307), .A2(rs2_val_gpr_w[23]), .ZN(n3491) );
  NAND2_X1 U3619 ( .A1(n3307), .A2(rs2_val_gpr_w[23]), .ZN(n3489) );
  OR2_X1 U3620 ( .A1(n3330), .A2(rs2_val_gpr_w[25]), .ZN(n3480) );
  NAND2_X1 U3621 ( .A1(n3330), .A2(rs2_val_gpr_w[25]), .ZN(n3478) );
  NOR2_X1 U3622 ( .A1(n3305), .A2(rs2_val_gpr_w[29]), .ZN(n3460) );
  NOR2_X1 U3623 ( .A1(n3347), .A2(rs2_val_gpr_w[30]), .ZN(n3465) );
  NAND2_X1 U3624 ( .A1(n3347), .A2(rs2_val_gpr_w[30]), .ZN(n3464) );
  NAND2_X1 U3625 ( .A1(n3342), .A2(rs1_val_gpr_w[29]), .ZN(n3469) );
  NAND2_X1 U3626 ( .A1(n3346), .A2(rs1_val_gpr_w[30]), .ZN(n3461) );
  AOI22_X1 U3627 ( .A1(alu_a_q[6]), .A2(alu_b_q[6]), .B1(n7165), .B2(n7164), 
        .ZN(n7187) );
  BUF_X2 U3628 ( .A(n5033), .Z(n3375) );
  INV_X1 U3629 ( .A(rs2_val_gpr_w[27]), .ZN(n3376) );
  BUF_X1 U3630 ( .A(rs1_val_gpr_w[7]), .Z(n3523) );
  OAI21_X1 U3631 ( .B1(n3812), .B2(n3781), .A(n7141), .ZN(n7164) );
  INV_X1 U3632 ( .A(rs2_val_gpr_w[9]), .ZN(n3377) );
  INV_X1 U3633 ( .A(rs2_val_gpr_w[14]), .ZN(n3378) );
  INV_X1 U3634 ( .A(rs1_val_gpr_w[6]), .ZN(n3379) );
  INV_X1 U3635 ( .A(rs1_val_gpr_w[1]), .ZN(n3380) );
  INV_X1 U3636 ( .A(rs2_val_gpr_w[10]), .ZN(n3381) );
  AND4_X1 U3637 ( .A1(n6050), .A2(n6049), .A3(n6048), .A4(n6047), .ZN(n3525)
         );
  INV_X1 U3638 ( .A(rs2_val_gpr_w[8]), .ZN(n3382) );
  INV_X1 U3639 ( .A(rs1_val_gpr_w[1]), .ZN(n3383) );
  INV_X1 U3640 ( .A(rs2_val_gpr_w[25]), .ZN(n3384) );
  INV_X1 U3641 ( .A(rs2_val_gpr_w[26]), .ZN(n3385) );
  INV_X1 U3642 ( .A(n7106), .ZN(n7119) );
  AND2_X2 U3643 ( .A1(n6790), .A2(n6813), .ZN(n6839) );
  AND2_X1 U3644 ( .A1(n5815), .A2(n5816), .ZN(n3411) );
  INV_X2 U3645 ( .A(n6492), .ZN(n6588) );
  INV_X1 U3646 ( .A(n7071), .ZN(n7072) );
  BUF_X1 U3647 ( .A(n5811), .Z(n4780) );
  AOI22_X1 U3648 ( .A1(n3286), .A2(reg_file[881]), .B1(n4806), .B2(
        reg_file[849]), .ZN(n6197) );
  OR2_X2 U3649 ( .A1(n3765), .A2(n7864), .ZN(n3842) );
  OR2_X2 U3650 ( .A1(n156), .A2(n7864), .ZN(n3764) );
  OAI22_X1 U3651 ( .A1(alu_a_q[1]), .A2(n3807), .B1(n7048), .B2(n7068), .ZN(
        n7071) );
  BUF_X1 U3652 ( .A(n3799), .Z(n4776) );
  BUF_X1 U3653 ( .A(n6385), .Z(n4802) );
  INV_X1 U3654 ( .A(n7990), .ZN(n7992) );
  NOR2_X1 U3655 ( .A1(n4942), .A2(mem_i_inst_i[16]), .ZN(n6384) );
  BUF_X1 U3656 ( .A(n6385), .Z(n4805) );
  NOR2_X1 U3657 ( .A1(alu_b_q[1]), .A2(n3779), .ZN(n7048) );
  NOR2_X1 U3658 ( .A1(n3774), .A2(n3808), .ZN(n7870) );
  NOR2_X1 U3659 ( .A1(n4945), .A2(n6604), .ZN(n6387) );
  INV_X1 U3660 ( .A(mem_i_inst_i[16]), .ZN(n6608) );
  INV_X1 U3661 ( .A(mem_i_inst_i[15]), .ZN(n6604) );
  INV_X1 U3662 ( .A(mem_i_inst_i[20]), .ZN(n6623) );
  INV_X1 U3663 ( .A(DP_OP_181_135_5161_n115), .ZN(n3434) );
  BUF_X1 U3664 ( .A(n7442), .Z(n4836) );
  BUF_X1 U3665 ( .A(n7642), .Z(n4840) );
  NOR3_X2 U3666 ( .A1(n3788), .A2(n3765), .A3(n154), .ZN(n7624) );
  OAI21_X2 U3667 ( .B1(n6958), .B2(n6957), .A(n3867), .ZN(n7012) );
  NOR2_X2 U3668 ( .A1(alu_b_q[3]), .A2(alu_b_q[2]), .ZN(n7414) );
  INV_X4 U3669 ( .A(n3796), .ZN(n4822) );
  INV_X1 U3670 ( .A(n3435), .ZN(n3391) );
  XNOR2_X1 U3671 ( .A(DP_OP_181_135_5161_n114), .B(n3391), .ZN(n3438) );
  XNOR2_X1 U3672 ( .A(DP_OP_181_135_5161_n116), .B(n3391), .ZN(n3447) );
  XNOR2_X1 U3673 ( .A(DP_OP_181_135_5161_n115), .B(n3391), .ZN(n3440) );
  AND2_X1 U3674 ( .A1(DP_OP_181_135_5161_n120), .A2(n3391), .ZN(n3484) );
  XNOR2_X1 U3675 ( .A(DP_OP_181_135_5161_n120), .B(n3391), .ZN(n3482) );
  NAND2_X1 U3676 ( .A1(DP_OP_181_135_5161_n117), .A2(n3391), .ZN(n3441) );
  NOR2_X1 U3677 ( .A1(DP_OP_181_135_5161_n117), .A2(n3391), .ZN(n3442) );
  INV_X1 U3678 ( .A(DP_OP_181_135_5161_n89), .ZN(n3435) );
  OAI21_X1 U3679 ( .B1(n6577), .B2(n4910), .A(n6560), .ZN(
        DP_OP_181_135_5161_n89) );
  NAND2_X1 U3680 ( .A1(DP_OP_181_135_5161_n24), .A2(n3396), .ZN(n3392) );
  NAND2_X1 U3681 ( .A1(n3393), .A2(n3392), .ZN(DP_OP_181_135_5161_n22) );
  AOI21_X1 U3682 ( .B1(n3415), .B2(n3398), .A(n3397), .ZN(n3463) );
  NOR3_X1 U3683 ( .A1(n3470), .A2(n3407), .A3(n3404), .ZN(n3400) );
  NOR2_X1 U3684 ( .A1(n3400), .A2(n3403), .ZN(n3402) );
  NAND2_X1 U3685 ( .A1(n3402), .A2(n3401), .ZN(n6456) );
  NAND2_X1 U3686 ( .A1(n3462), .A2(n3461), .ZN(n3409) );
  NAND2_X1 U3687 ( .A1(n3461), .A2(n3469), .ZN(n3410) );
  NAND2_X1 U3688 ( .A1(sub_x_59_n7), .A2(n3414), .ZN(n3412) );
  NAND2_X1 U3689 ( .A1(n3412), .A2(n3413), .ZN(n3472) );
  NAND2_X1 U3690 ( .A1(n3479), .A2(n3478), .ZN(n3425) );
  OAI21_X1 U3691 ( .B1(n3427), .B2(n3509), .A(n3426), .ZN(n3501) );
  OR2_X1 U3692 ( .A1(n3310), .A2(rs1_val_gpr_w[23]), .ZN(n3426) );
  AOI21_X1 U3693 ( .B1(n3502), .B2(n3573), .A(n3510), .ZN(n3427) );
  AND2_X1 U3694 ( .A1(DP_OP_181_135_5161_n107), .A2(DP_OP_181_135_5161_n86), 
        .ZN(n3431) );
  NAND2_X1 U3695 ( .A1(sub_x_60_n8), .A2(n3480), .ZN(n3479) );
  INV_X1 U3696 ( .A(n3436), .ZN(DP_OP_181_135_5161_n8) );
  AOI22_X1 U3697 ( .A1(DP_OP_181_135_5161_n9), .A2(n3437), .B1(n3391), .B2(
        DP_OP_181_135_5161_n114), .ZN(n3436) );
  NOR2_X1 U3698 ( .A1(DP_OP_181_135_5161_n115), .A2(n3391), .ZN(n3439) );
  AND2_X1 U3699 ( .A1(DP_OP_181_135_5161_n116), .A2(n3391), .ZN(n3445) );
  OAI21_X1 U3700 ( .B1(n3449), .B2(n3450), .A(n3448), .ZN(
        DP_OP_181_135_5161_n30) );
  NAND2_X1 U3701 ( .A1(DP_OP_181_135_5161_n92), .A2(C1_Z_2), .ZN(n3448) );
  NOR2_X1 U3702 ( .A1(DP_OP_181_135_5161_n92), .A2(C1_Z_2), .ZN(n3449) );
  AOI21_X1 U3703 ( .B1(n3452), .B2(DP_OP_181_135_5161_n32), .A(n3451), .ZN(
        n3450) );
  NAND3_X1 U3704 ( .A1(n3454), .A2(n6476), .A3(n3453), .ZN(n2885) );
  AND2_X1 U3705 ( .A1(DP_OP_181_135_5161_n95), .A2(DP_OP_181_135_5161_n74), 
        .ZN(n3458) );
  NAND2_X1 U3706 ( .A1(n3472), .A2(n3471), .ZN(n3470) );
  XNOR2_X1 U3707 ( .A(n3463), .B(sub_x_60_n1), .ZN(u_branch_N120) );
  OAI21_X1 U3708 ( .B1(n3468), .B2(n3467), .A(n3466), .ZN(sub_x_59_n8) );
  NAND2_X1 U3709 ( .A1(n3336), .A2(rs1_val_gpr_w[24]), .ZN(n3466) );
  NOR2_X1 U3710 ( .A1(n3336), .A2(rs1_val_gpr_w[24]), .ZN(n3467) );
  NAND2_X1 U3711 ( .A1(n3473), .A2(n3491), .ZN(n3490) );
  NAND2_X1 U3712 ( .A1(n3475), .A2(n3474), .ZN(n3473) );
  NAND2_X1 U3713 ( .A1(n3344), .A2(rs2_val_gpr_w[22]), .ZN(n3474) );
  NAND2_X1 U3714 ( .A1(sub_x_60_n11), .A2(n3476), .ZN(n3475) );
  OR2_X1 U3715 ( .A1(n3344), .A2(rs2_val_gpr_w[22]), .ZN(n3476) );
  NAND2_X1 U3716 ( .A1(n3490), .A2(n3489), .ZN(sub_x_60_n9) );
  NAND2_X1 U3717 ( .A1(sub_x_59_n8), .A2(n3499), .ZN(n3498) );
  NAND2_X1 U3718 ( .A1(n3498), .A2(n3497), .ZN(sub_x_59_n7) );
  NAND2_X1 U3719 ( .A1(n3493), .A2(n3492), .ZN(DP_OP_181_135_5161_n29) );
  NAND2_X1 U3720 ( .A1(DP_OP_181_135_5161_n30), .A2(n3494), .ZN(n3493) );
  NAND2_X1 U3721 ( .A1(n3495), .A2(n6580), .ZN(n3494) );
  INV_X1 U3722 ( .A(DP_OP_181_135_5161_n93), .ZN(n3495) );
  AOI21_X1 U3723 ( .B1(n3503), .B2(n3527), .A(n3507), .ZN(n3506) );
  AOI21_X1 U3724 ( .B1(n3508), .B2(n3506), .A(n3504), .ZN(sub_x_60_n11) );
  NOR2_X1 U3725 ( .A1(sub_x_60_n12), .A2(n3505), .ZN(n3504) );
  INV_X1 U3726 ( .A(n3723), .ZN(n3505) );
  NAND2_X1 U3727 ( .A1(n3723), .A2(n3540), .ZN(n3507) );
  AOI21_X1 U3728 ( .B1(n3514), .B2(n3513), .A(n3512), .ZN(n3511) );
  INV_X1 U3729 ( .A(n3515), .ZN(n3514) );
  OAI21_X1 U3730 ( .B1(sub_x_59_n28), .B2(n3578), .A(sub_x_59_n29), .ZN(n3515)
         );
  BUF_X1 U3731 ( .A(n5809), .Z(n3519) );
  INV_X1 U3732 ( .A(mem_i_inst_i[17]), .ZN(n3520) );
  NAND4_X1 U3733 ( .A1(n4969), .A2(n4968), .A3(n4967), .A4(n4966), .ZN(
        rs1_val_gpr_w[0]) );
  INV_X1 U3734 ( .A(n3317), .ZN(n3522) );
  INV_X1 U3735 ( .A(n3317), .ZN(n4813) );
  INV_X1 U3736 ( .A(n3288), .ZN(n3524) );
  AND4_X1 U3737 ( .A1(n4969), .A2(n4968), .A3(n4967), .A4(n4966), .ZN(n3526)
         );
  AOI21_X1 U3738 ( .B1(n6456), .B2(n6741), .A(n6455), .ZN(n6459) );
  NOR2_X1 U3739 ( .A1(n6459), .A2(n4719), .ZN(n4718) );
  OR2_X1 U3740 ( .A1(n6454), .A2(n4713), .ZN(n4712) );
  NOR2_X1 U3741 ( .A1(rs2_val_gpr_w[1]), .A2(n3383), .ZN(sub_x_60_n92) );
  NAND2_X1 U3742 ( .A1(rs2_val_gpr_w[1]), .A2(n3383), .ZN(sub_x_60_n93) );
  NOR2_X1 U3743 ( .A1(rs2_val_gpr_w[0]), .A2(n3526), .ZN(sub_x_60_n94) );
  AND2_X1 U3744 ( .A1(n3543), .A2(n3556), .ZN(n3535) );
  INV_X1 U3745 ( .A(n3535), .ZN(n3536) );
  AND2_X1 U3746 ( .A1(rs2_val_gpr_w[16]), .A2(n3339), .ZN(n3541) );
  OR2_X1 U3747 ( .A1(rs2_val_gpr_w[10]), .A2(n3525), .ZN(n3543) );
  AND2_X1 U3748 ( .A1(rs2_val_gpr_w[15]), .A2(n3304), .ZN(n3545) );
  AND2_X1 U3749 ( .A1(rs2_val_gpr_w[7]), .A2(n3327), .ZN(n3546) );
  OR2_X1 U3750 ( .A1(rs2_val_gpr_w[2]), .A2(n3329), .ZN(n3547) );
  OR2_X1 U3751 ( .A1(rs2_val_gpr_w[4]), .A2(n3324), .ZN(n3548) );
  OR2_X1 U3752 ( .A1(rs2_val_gpr_w[18]), .A2(n3334), .ZN(n3550) );
  AND2_X1 U3753 ( .A1(rs2_val_gpr_w[2]), .A2(n3329), .ZN(n3551) );
  AND2_X1 U3754 ( .A1(rs2_val_gpr_w[6]), .A2(n3379), .ZN(n3552) );
  AND2_X1 U3755 ( .A1(rs2_val_gpr_w[4]), .A2(n3324), .ZN(n3553) );
  OR2_X1 U3756 ( .A1(rs2_val_gpr_w[15]), .A2(n3304), .ZN(n3555) );
  OR2_X1 U3757 ( .A1(rs2_val_gpr_w[11]), .A2(n3289), .ZN(n3556) );
  OR2_X1 U3758 ( .A1(rs2_val_gpr_w[13]), .A2(n3290), .ZN(n3557) );
  OR2_X1 U3759 ( .A1(rs2_val_gpr_w[7]), .A2(n3327), .ZN(n3558) );
  AOI21_X1 U3760 ( .B1(n3552), .B2(n3558), .A(n3546), .ZN(n3531) );
  OAI21_X1 U3761 ( .B1(sub_x_60_n92), .B2(sub_x_60_n94), .A(sub_x_60_n93), 
        .ZN(n3532) );
  AOI21_X1 U3762 ( .B1(n3547), .B2(n3532), .A(n3551), .ZN(n3533) );
  OAI21_X1 U3763 ( .B1(n3533), .B2(sub_x_60_n84), .A(n3691), .ZN(n3534) );
  AOI21_X1 U3764 ( .B1(n3534), .B2(n3548), .A(n3553), .ZN(sub_x_60_n78) );
  INV_X1 U3765 ( .A(sub_x_59_n41), .ZN(sub_x_59_n39) );
  INV_X1 U3766 ( .A(sub_x_59_n65), .ZN(sub_x_59_n63) );
  NOR2_X1 U3767 ( .A1(n3302), .A2(rs1_val_gpr_w[1]), .ZN(sub_x_59_n92) );
  NAND2_X1 U3768 ( .A1(n3302), .A2(rs1_val_gpr_w[1]), .ZN(sub_x_59_n93) );
  NAND2_X1 U3769 ( .A1(n3568), .A2(n3567), .ZN(sub_x_59_n59) );
  NAND3_X1 U3770 ( .A1(n3564), .A2(n3598), .A3(n3580), .ZN(n3568) );
  NAND2_X1 U3771 ( .A1(n3571), .A2(n3570), .ZN(n3559) );
  NAND3_X1 U3772 ( .A1(sub_x_59_n59), .A2(n3600), .A3(n3579), .ZN(n3571) );
  AND2_X1 U3773 ( .A1(n3312), .A2(rs1_val_gpr_w[21]), .ZN(n3577) );
  AND3_X1 U3774 ( .A1(n3583), .A2(n3597), .A3(sub_x_59_n39), .ZN(n3579) );
  AND3_X1 U3775 ( .A1(n3596), .A2(n3592), .A3(sub_x_59_n63), .ZN(n3580) );
  AND2_X1 U3776 ( .A1(n3377), .A2(rs1_val_gpr_w[9]), .ZN(n3585) );
  AND2_X1 U3777 ( .A1(n3322), .A2(rs1_val_gpr_w[11]), .ZN(n3586) );
  AND2_X1 U3778 ( .A1(n3311), .A2(rs1_val_gpr_w[15]), .ZN(n3587) );
  AND2_X1 U3779 ( .A1(n3292), .A2(rs1_val_gpr_w[7]), .ZN(n3588) );
  AND2_X1 U3780 ( .A1(n3291), .A2(rs1_val_gpr_w[13]), .ZN(n3589) );
  AND2_X1 U3781 ( .A1(n3309), .A2(rs1_val_gpr_w[2]), .ZN(n3590) );
  OR2_X1 U3782 ( .A1(n3325), .A2(rs1_val_gpr_w[4]), .ZN(n3591) );
  OR2_X1 U3783 ( .A1(n3313), .A2(rs1_val_gpr_w[6]), .ZN(n3592) );
  OR2_X1 U3784 ( .A1(n3350), .A2(rs1_val_gpr_w[12]), .ZN(n3593) );
  OR2_X1 U3785 ( .A1(n3332), .A2(rs1_val_gpr_w[19]), .ZN(n3594) );
  OR2_X1 U3786 ( .A1(n3312), .A2(rs1_val_gpr_w[21]), .ZN(n3595) );
  OR2_X1 U3787 ( .A1(n3292), .A2(rs1_val_gpr_w[7]), .ZN(n3596) );
  OR2_X1 U3788 ( .A1(n3291), .A2(rs1_val_gpr_w[13]), .ZN(n3597) );
  OR2_X1 U3789 ( .A1(n3377), .A2(rs1_val_gpr_w[9]), .ZN(n3598) );
  OR2_X1 U3790 ( .A1(n3322), .A2(rs1_val_gpr_w[11]), .ZN(n3599) );
  OR2_X1 U3791 ( .A1(n3311), .A2(rs1_val_gpr_w[15]), .ZN(n3600) );
  AND2_X1 U3792 ( .A1(n3325), .A2(rs1_val_gpr_w[4]), .ZN(n3601) );
  OR2_X1 U3793 ( .A1(n3309), .A2(rs1_val_gpr_w[2]), .ZN(n3602) );
  AND2_X1 U3794 ( .A1(n3381), .A2(rs1_val_gpr_w[10]), .ZN(n3603) );
  AND2_X1 U3795 ( .A1(n3313), .A2(rs1_val_gpr_w[6]), .ZN(n3604) );
  OAI21_X1 U3796 ( .B1(sub_x_59_n94), .B2(sub_x_59_n92), .A(sub_x_59_n93), 
        .ZN(n3574) );
  AOI21_X1 U3797 ( .B1(n3574), .B2(n3602), .A(n3590), .ZN(n3575) );
  OAI21_X1 U3798 ( .B1(n3575), .B2(sub_x_59_n84), .A(sub_x_59_n85), .ZN(n3576)
         );
  AOI21_X1 U3799 ( .B1(n3576), .B2(n3591), .A(n3601), .ZN(sub_x_59_n78) );
  OAI21_X1 U3800 ( .B1(sub_x_59_n78), .B2(sub_x_59_n76), .A(sub_x_59_n77), 
        .ZN(n3564) );
  AOI21_X1 U3801 ( .B1(n3604), .B2(n3596), .A(n3588), .ZN(n3565) );
  OAI21_X1 U3802 ( .B1(n3565), .B2(sub_x_59_n65), .A(n3582), .ZN(n3566) );
  AOI21_X1 U3803 ( .B1(n3566), .B2(n3598), .A(n3585), .ZN(n3567) );
  AOI21_X1 U3804 ( .B1(n3603), .B2(n3599), .A(n3586), .ZN(n3560) );
  INV_X1 U3805 ( .A(n3593), .ZN(n3561) );
  OAI21_X1 U3806 ( .B1(n3560), .B2(n3561), .A(n3584), .ZN(n3562) );
  AOI21_X1 U3807 ( .B1(n3562), .B2(n3597), .A(n3589), .ZN(n3563) );
  OAI21_X1 U3808 ( .B1(n3563), .B2(sub_x_59_n41), .A(n3581), .ZN(n3569) );
  AOI21_X1 U3809 ( .B1(n3569), .B2(n3600), .A(n3587), .ZN(n3570) );
  AOI21_X1 U3810 ( .B1(n3572), .B2(n3595), .A(n3577), .ZN(n3573) );
  NOR2_X1 U3811 ( .A1(rs2_val_gpr_w[29]), .A2(n3305), .ZN(n3606) );
  NAND2_X1 U3812 ( .A1(rs1_val_gpr_w[31]), .A2(n3298), .ZN(n3605) );
  OAI21_X1 U3813 ( .B1(rs2_val_gpr_w[30]), .B2(n3347), .A(n3605), .ZN(n3660)
         );
  AOI211_X1 U3814 ( .C1(rs1_val_gpr_w[28]), .C2(n3348), .A(n3606), .B(n3660), 
        .ZN(n3666) );
  NOR2_X1 U3815 ( .A1(rs2_val_gpr_w[25]), .A2(n3330), .ZN(n3664) );
  NOR2_X1 U3816 ( .A1(n3331), .A2(rs2_val_gpr_w[27]), .ZN(n3662) );
  AOI21_X1 U3817 ( .B1(n3385), .B2(rs1_val_gpr_w[26]), .A(n3662), .ZN(n3607)
         );
  AOI211_X1 U3818 ( .C1(rs1_val_gpr_w[24]), .C2(n3336), .A(n3664), .B(n3679), 
        .ZN(n3608) );
  NAND2_X1 U3819 ( .A1(n3666), .A2(n3608), .ZN(n3676) );
  NOR2_X1 U3820 ( .A1(rs2_val_gpr_w[9]), .A2(n3308), .ZN(n3629) );
  NOR2_X1 U3821 ( .A1(rs2_val_gpr_w[11]), .A2(n3289), .ZN(n3627) );
  AOI21_X1 U3822 ( .B1(n3381), .B2(rs1_val_gpr_w[10]), .A(n3627), .ZN(n3609)
         );
  NOR2_X1 U3823 ( .A1(rs2_val_gpr_w[8]), .A2(n3321), .ZN(n3612) );
  NOR2_X1 U3824 ( .A1(rs2_val_gpr_w[15]), .A2(n3304), .ZN(n3610) );
  AOI21_X1 U3825 ( .B1(rs1_val_gpr_w[14]), .B2(n3378), .A(n3610), .ZN(n3638)
         );
  NAND2_X1 U3826 ( .A1(rs1_val_gpr_w[13]), .A2(n3291), .ZN(n3611) );
  OAI211_X1 U3827 ( .C1(rs2_val_gpr_w[12]), .C2(n3351), .A(n3638), .B(n3611), 
        .ZN(n3631) );
  OR4_X1 U3828 ( .A1(n3629), .A2(n3677), .A3(n3612), .A4(n3631), .ZN(n3641) );
  OAI21_X1 U3829 ( .B1(rs2_val_gpr_w[5]), .B2(n3306), .A(rs2_val_gpr_w[4]), 
        .ZN(n3613) );
  OAI22_X1 U3830 ( .A1(rs1_val_gpr_w[4]), .A2(n3613), .B1(rs1_val_gpr_w[5]), 
        .B2(n3303), .ZN(n3625) );
  NOR2_X1 U3831 ( .A1(rs2_val_gpr_w[7]), .A2(n3327), .ZN(n3614) );
  AOI21_X1 U3832 ( .B1(rs1_val_gpr_w[6]), .B2(n3313), .A(n3614), .ZN(n3624) );
  OAI21_X1 U3833 ( .B1(rs2_val_gpr_w[3]), .B2(n3288), .A(rs2_val_gpr_w[2]), 
        .ZN(n3618) );
  OAI21_X1 U3834 ( .B1(rs2_val_gpr_w[1]), .B2(n3380), .A(rs2_val_gpr_w[0]), 
        .ZN(n3615) );
  OAI22_X1 U3835 ( .A1(n3521), .A2(n3615), .B1(rs1_val_gpr_w[1]), .B2(n3302), 
        .ZN(n3616) );
  OAI221_X1 U3836 ( .B1(rs2_val_gpr_w[3]), .B2(n3288), .C1(rs2_val_gpr_w[2]), 
        .C2(n3329), .A(n3616), .ZN(n3617) );
  OAI221_X1 U3837 ( .B1(rs1_val_gpr_w[3]), .B2(n3299), .C1(rs1_val_gpr_w[2]), 
        .C2(n3618), .A(n3617), .ZN(n3619) );
  OAI21_X1 U3838 ( .B1(rs2_val_gpr_w[5]), .B2(n3306), .A(n3619), .ZN(n3620) );
  AOI21_X1 U3839 ( .B1(rs1_val_gpr_w[4]), .B2(n3325), .A(n3620), .ZN(n3623) );
  OAI21_X1 U3840 ( .B1(rs2_val_gpr_w[7]), .B2(n3327), .A(rs2_val_gpr_w[6]), 
        .ZN(n3621) );
  OAI22_X1 U3841 ( .A1(rs1_val_gpr_w[6]), .A2(n3621), .B1(n3523), .B2(n3292), 
        .ZN(n3622) );
  AOI221_X1 U3842 ( .B1(n3625), .B2(n3624), .C1(n3623), .C2(n3624), .A(n3622), 
        .ZN(n3640) );
  OAI21_X1 U3843 ( .B1(rs2_val_gpr_w[13]), .B2(n3290), .A(rs2_val_gpr_w[12]), 
        .ZN(n3626) );
  OAI22_X1 U3844 ( .A1(rs1_val_gpr_w[12]), .A2(n3626), .B1(rs1_val_gpr_w[13]), 
        .B2(n3291), .ZN(n3637) );
  NOR2_X1 U3845 ( .A1(n3627), .A2(rs1_val_gpr_w[10]), .ZN(n3628) );
  AOI22_X1 U3846 ( .A1(rs2_val_gpr_w[11]), .A2(n3289), .B1(rs2_val_gpr_w[10]), 
        .B2(n3628), .ZN(n3633) );
  NOR2_X1 U3847 ( .A1(n3629), .A2(rs1_val_gpr_w[8]), .ZN(n3630) );
  AOI22_X1 U3848 ( .A1(n3630), .A2(rs2_val_gpr_w[8]), .B1(rs2_val_gpr_w[9]), 
        .B2(n3308), .ZN(n3632) );
  AOI221_X1 U3849 ( .B1(n3677), .B2(n3633), .C1(n3632), .C2(n3633), .A(n3631), 
        .ZN(n3636) );
  OAI21_X1 U3850 ( .B1(rs2_val_gpr_w[15]), .B2(n3304), .A(rs2_val_gpr_w[14]), 
        .ZN(n3634) );
  OAI22_X1 U3851 ( .A1(rs1_val_gpr_w[14]), .A2(n3634), .B1(rs1_val_gpr_w[15]), 
        .B2(n3311), .ZN(n3635) );
  AOI211_X1 U3852 ( .C1(n3638), .C2(n3637), .A(n3636), .B(n3635), .ZN(n3639)
         );
  OAI21_X1 U3853 ( .B1(n3641), .B2(n3640), .A(n3639), .ZN(n3646) );
  NOR2_X1 U3854 ( .A1(rs2_val_gpr_w[17]), .A2(n3300), .ZN(n3650) );
  NOR2_X1 U3855 ( .A1(rs2_val_gpr_w[23]), .A2(n3307), .ZN(n3642) );
  AOI21_X1 U3856 ( .B1(rs1_val_gpr_w[22]), .B2(n3343), .A(n3642), .ZN(n3659)
         );
  NAND2_X1 U3857 ( .A1(rs1_val_gpr_w[21]), .A2(n3312), .ZN(n3643) );
  OAI211_X1 U3858 ( .C1(rs2_val_gpr_w[20]), .C2(n3341), .A(n3659), .B(n3643), 
        .ZN(n3652) );
  NOR2_X1 U3859 ( .A1(rs2_val_gpr_w[19]), .A2(n3349), .ZN(n3648) );
  AOI21_X1 U3860 ( .B1(n3337), .B2(rs1_val_gpr_w[18]), .A(n3648), .ZN(n3644)
         );
  AOI211_X1 U3861 ( .C1(rs1_val_gpr_w[16]), .C2(n3338), .A(n3652), .B(n3678), 
        .ZN(n3645) );
  NAND3_X1 U3862 ( .A1(n3646), .A2(sub_x_60_n28), .A3(n3645), .ZN(n3675) );
  OAI21_X1 U3863 ( .B1(rs2_val_gpr_w[21]), .B2(n3301), .A(rs2_val_gpr_w[20]), 
        .ZN(n3647) );
  OAI22_X1 U3864 ( .A1(rs1_val_gpr_w[20]), .A2(n3647), .B1(rs1_val_gpr_w[21]), 
        .B2(n3312), .ZN(n3658) );
  NOR2_X1 U3865 ( .A1(rs1_val_gpr_w[18]), .A2(n3648), .ZN(n3649) );
  AOI22_X1 U3866 ( .A1(rs2_val_gpr_w[18]), .A2(n3649), .B1(rs2_val_gpr_w[19]), 
        .B2(n3349), .ZN(n3654) );
  NOR2_X1 U3867 ( .A1(rs1_val_gpr_w[16]), .A2(n3650), .ZN(n3651) );
  AOI22_X1 U3868 ( .A1(rs2_val_gpr_w[16]), .A2(n3651), .B1(rs2_val_gpr_w[17]), 
        .B2(n3300), .ZN(n3653) );
  AOI221_X1 U3869 ( .B1(n3678), .B2(n3654), .C1(n3653), .C2(n3654), .A(n3652), 
        .ZN(n3657) );
  OAI21_X1 U3870 ( .B1(rs2_val_gpr_w[23]), .B2(n3307), .A(rs2_val_gpr_w[22]), 
        .ZN(n3655) );
  OAI22_X1 U3871 ( .A1(rs1_val_gpr_w[22]), .A2(n3655), .B1(rs1_val_gpr_w[23]), 
        .B2(n3310), .ZN(n3656) );
  AOI211_X1 U3872 ( .C1(n3659), .C2(n3658), .A(n3657), .B(n3656), .ZN(n3674)
         );
  OAI21_X1 U3873 ( .B1(rs2_val_gpr_w[29]), .B2(n3305), .A(rs2_val_gpr_w[28]), 
        .ZN(n3661) );
  OAI22_X1 U3874 ( .A1(rs1_val_gpr_w[28]), .A2(n3661), .B1(rs1_val_gpr_w[29]), 
        .B2(n3342), .ZN(n3672) );
  NOR2_X1 U3875 ( .A1(rs1_val_gpr_w[26]), .A2(n3662), .ZN(n3663) );
  AOI22_X1 U3876 ( .A1(rs2_val_gpr_w[26]), .A2(n3663), .B1(rs2_val_gpr_w[27]), 
        .B2(n3331), .ZN(n3668) );
  NOR2_X1 U3877 ( .A1(rs1_val_gpr_w[24]), .A2(n3664), .ZN(n3665) );
  AOI22_X1 U3878 ( .A1(rs2_val_gpr_w[24]), .A2(n3665), .B1(rs2_val_gpr_w[25]), 
        .B2(n3330), .ZN(n3667) );
  AOI221_X1 U3879 ( .B1(n3679), .B2(n3668), .C1(n3667), .C2(n3668), .A(n3681), 
        .ZN(n3671) );
  OAI21_X1 U3880 ( .B1(rs2_val_gpr_w[31]), .B2(n3345), .A(rs2_val_gpr_w[30]), 
        .ZN(n3669) );
  OAI22_X1 U3881 ( .A1(rs1_val_gpr_w[30]), .A2(n3669), .B1(rs1_val_gpr_w[31]), 
        .B2(n3298), .ZN(n3670) );
  AOI211_X1 U3882 ( .C1(n3680), .C2(n3672), .A(n3671), .B(n3670), .ZN(n3673)
         );
  OAI221_X1 U3883 ( .B1(n3676), .B2(n3675), .C1(n3676), .C2(n3674), .A(n3673), 
        .ZN(u_branch_N125) );
  INV_X1 U3884 ( .A(n3607), .ZN(n3679) );
  INV_X1 U3885 ( .A(n3609), .ZN(n3677) );
  INV_X1 U3886 ( .A(n3644), .ZN(n3678) );
  INV_X1 U3887 ( .A(n3660), .ZN(n3680) );
  INV_X1 U3888 ( .A(n3666), .ZN(n3681) );
  NOR2_X1 U3889 ( .A1(rs1_val_gpr_w[29]), .A2(n3342), .ZN(n3683) );
  NAND2_X1 U3890 ( .A1(rs2_val_gpr_w[31]), .A2(n3345), .ZN(n3682) );
  OAI21_X1 U3891 ( .B1(rs1_val_gpr_w[30]), .B2(n3346), .A(n3682), .ZN(n3740)
         );
  AOI211_X1 U3892 ( .C1(rs2_val_gpr_w[28]), .C2(n3320), .A(n3683), .B(n3740), 
        .ZN(n3746) );
  NOR2_X1 U3893 ( .A1(rs1_val_gpr_w[25]), .A2(n3384), .ZN(n3744) );
  NOR2_X1 U3894 ( .A1(n3376), .A2(rs1_val_gpr_w[27]), .ZN(n3742) );
  AOI21_X1 U3895 ( .B1(n3333), .B2(rs2_val_gpr_w[26]), .A(n3742), .ZN(n3684)
         );
  AOI211_X1 U3896 ( .C1(rs2_val_gpr_w[24]), .C2(n3335), .A(n3744), .B(n3759), 
        .ZN(n3685) );
  NAND2_X1 U3897 ( .A1(n3746), .A2(n3685), .ZN(n3756) );
  NAND2_X1 U3898 ( .A1(rs2_val_gpr_w[7]), .A2(n3327), .ZN(n3687) );
  NAND3_X1 U3899 ( .A1(n3313), .A2(n3687), .A3(rs1_val_gpr_w[6]), .ZN(n3686)
         );
  OAI21_X1 U3900 ( .B1(rs2_val_gpr_w[7]), .B2(n3327), .A(n3686), .ZN(n3706) );
  OAI21_X1 U3901 ( .B1(rs1_val_gpr_w[6]), .B2(n3313), .A(n3687), .ZN(n3699) );
  NOR2_X1 U3902 ( .A1(rs1_val_gpr_w[5]), .A2(n3303), .ZN(n3689) );
  NOR2_X1 U3903 ( .A1(n3689), .A2(rs2_val_gpr_w[4]), .ZN(n3688) );
  AOI22_X1 U3904 ( .A1(n3688), .A2(rs1_val_gpr_w[4]), .B1(rs1_val_gpr_w[5]), 
        .B2(n3303), .ZN(n3698) );
  AOI21_X1 U3905 ( .B1(rs2_val_gpr_w[4]), .B2(n3324), .A(n3689), .ZN(n3696) );
  OAI21_X1 U3906 ( .B1(rs2_val_gpr_w[1]), .B2(n3383), .A(rs2_val_gpr_w[0]), 
        .ZN(n3690) );
  OAI22_X1 U3907 ( .A1(n3521), .A2(n3690), .B1(rs1_val_gpr_w[1]), .B2(n3302), 
        .ZN(n3694) );
  NAND2_X1 U3908 ( .A1(rs2_val_gpr_w[3]), .A2(n3288), .ZN(n3691) );
  OAI21_X1 U3909 ( .B1(rs1_val_gpr_w[2]), .B2(n3309), .A(n3691), .ZN(n3693) );
  NAND3_X1 U3910 ( .A1(n3691), .A2(n3309), .A3(rs1_val_gpr_w[2]), .ZN(n3692)
         );
  OAI221_X1 U3911 ( .B1(rs2_val_gpr_w[3]), .B2(n3288), .C1(n3694), .C2(n3693), 
        .A(n3692), .ZN(n3695) );
  NAND2_X1 U3912 ( .A1(n3696), .A2(n3695), .ZN(n3697) );
  OAI22_X1 U3913 ( .A1(n3699), .A2(n3698), .B1(n3699), .B2(n3697), .ZN(n3705)
         );
  NOR2_X1 U3914 ( .A1(rs1_val_gpr_w[15]), .A2(n3311), .ZN(n3700) );
  AOI21_X1 U3915 ( .B1(rs2_val_gpr_w[14]), .B2(n3323), .A(n3700), .ZN(n3719)
         );
  NAND2_X1 U3916 ( .A1(rs2_val_gpr_w[13]), .A2(n3290), .ZN(n3701) );
  OAI211_X1 U3917 ( .C1(rs1_val_gpr_w[12]), .C2(n3350), .A(n3719), .B(n3701), 
        .ZN(n3712) );
  NOR2_X1 U3918 ( .A1(rs1_val_gpr_w[8]), .A2(n3382), .ZN(n3703) );
  NOR2_X1 U3919 ( .A1(rs1_val_gpr_w[9]), .A2(n3377), .ZN(n3710) );
  NOR2_X1 U3920 ( .A1(rs1_val_gpr_w[11]), .A2(n3322), .ZN(n3708) );
  AOI21_X1 U3921 ( .B1(n3525), .B2(rs2_val_gpr_w[10]), .A(n3708), .ZN(n3702)
         );
  NOR4_X1 U3922 ( .A1(n3712), .A2(n3703), .A3(n3710), .A4(n3757), .ZN(n3704)
         );
  OAI21_X1 U3923 ( .B1(n3706), .B2(n3705), .A(n3704), .ZN(n3721) );
  OAI21_X1 U3924 ( .B1(rs1_val_gpr_w[13]), .B2(n3291), .A(rs1_val_gpr_w[12]), 
        .ZN(n3707) );
  OAI22_X1 U3925 ( .A1(rs2_val_gpr_w[12]), .A2(n3707), .B1(n3290), .B2(
        rs2_val_gpr_w[13]), .ZN(n3718) );
  NOR2_X1 U3926 ( .A1(rs2_val_gpr_w[10]), .A2(n3708), .ZN(n3709) );
  AOI22_X1 U3927 ( .A1(rs1_val_gpr_w[10]), .A2(n3709), .B1(rs1_val_gpr_w[11]), 
        .B2(n3322), .ZN(n3714) );
  NOR2_X1 U3928 ( .A1(rs2_val_gpr_w[8]), .A2(n3710), .ZN(n3711) );
  AOI22_X1 U3929 ( .A1(rs1_val_gpr_w[8]), .A2(n3711), .B1(rs1_val_gpr_w[9]), 
        .B2(n3377), .ZN(n3713) );
  AOI221_X1 U3930 ( .B1(n3757), .B2(n3714), .C1(n3713), .C2(n3714), .A(n3712), 
        .ZN(n3717) );
  OAI21_X1 U3931 ( .B1(rs1_val_gpr_w[15]), .B2(n3311), .A(rs1_val_gpr_w[14]), 
        .ZN(n3715) );
  OAI22_X1 U3932 ( .A1(rs2_val_gpr_w[14]), .A2(n3715), .B1(rs2_val_gpr_w[15]), 
        .B2(n3304), .ZN(n3716) );
  AOI211_X1 U3933 ( .C1(n3719), .C2(n3718), .A(n3717), .B(n3716), .ZN(n3720)
         );
  NOR2_X1 U3934 ( .A1(rs1_val_gpr_w[17]), .A2(n3340), .ZN(n3730) );
  AOI21_X1 U3935 ( .B1(n3721), .B2(n3720), .A(n3730), .ZN(n3726) );
  NOR2_X1 U3936 ( .A1(rs1_val_gpr_w[23]), .A2(n3310), .ZN(n3722) );
  AOI21_X1 U3937 ( .B1(rs2_val_gpr_w[22]), .B2(n3344), .A(n3722), .ZN(n3739)
         );
  NAND2_X1 U3938 ( .A1(rs2_val_gpr_w[21]), .A2(n3301), .ZN(n3723) );
  OAI211_X1 U3939 ( .C1(rs1_val_gpr_w[20]), .C2(n3326), .A(n3739), .B(n3723), 
        .ZN(n3732) );
  NOR2_X1 U3940 ( .A1(rs1_val_gpr_w[19]), .A2(n3332), .ZN(n3728) );
  AOI21_X1 U3941 ( .B1(n3334), .B2(rs2_val_gpr_w[18]), .A(n3728), .ZN(n3724)
         );
  AOI211_X1 U3942 ( .C1(rs2_val_gpr_w[16]), .C2(n3339), .A(n3732), .B(n3758), 
        .ZN(n3725) );
  NAND2_X1 U3943 ( .A1(n3726), .A2(n3725), .ZN(n3755) );
  OAI21_X1 U3944 ( .B1(rs1_val_gpr_w[21]), .B2(n3312), .A(rs1_val_gpr_w[20]), 
        .ZN(n3727) );
  OAI22_X1 U3945 ( .A1(rs2_val_gpr_w[20]), .A2(n3727), .B1(rs2_val_gpr_w[21]), 
        .B2(n3301), .ZN(n3738) );
  NOR2_X1 U3946 ( .A1(rs2_val_gpr_w[18]), .A2(n3728), .ZN(n3729) );
  AOI22_X1 U3947 ( .A1(rs1_val_gpr_w[18]), .A2(n3729), .B1(rs1_val_gpr_w[19]), 
        .B2(n3332), .ZN(n3734) );
  NOR2_X1 U3948 ( .A1(rs2_val_gpr_w[16]), .A2(n3730), .ZN(n3731) );
  AOI22_X1 U3949 ( .A1(rs1_val_gpr_w[16]), .A2(n3731), .B1(rs1_val_gpr_w[17]), 
        .B2(n3340), .ZN(n3733) );
  AOI221_X1 U3950 ( .B1(n3758), .B2(n3734), .C1(n3733), .C2(n3734), .A(n3732), 
        .ZN(n3737) );
  OAI21_X1 U3951 ( .B1(rs1_val_gpr_w[23]), .B2(n3310), .A(rs1_val_gpr_w[22]), 
        .ZN(n3735) );
  OAI22_X1 U3952 ( .A1(rs2_val_gpr_w[22]), .A2(n3735), .B1(rs2_val_gpr_w[23]), 
        .B2(n3307), .ZN(n3736) );
  AOI211_X1 U3953 ( .C1(n3739), .C2(n3738), .A(n3737), .B(n3736), .ZN(n3754)
         );
  OAI21_X1 U3954 ( .B1(rs1_val_gpr_w[29]), .B2(n3342), .A(rs1_val_gpr_w[28]), 
        .ZN(n3741) );
  OAI22_X1 U3955 ( .A1(rs2_val_gpr_w[28]), .A2(n3741), .B1(rs2_val_gpr_w[29]), 
        .B2(n3305), .ZN(n3752) );
  NOR2_X1 U3956 ( .A1(rs2_val_gpr_w[26]), .A2(n3742), .ZN(n3743) );
  AOI22_X1 U3957 ( .A1(rs1_val_gpr_w[26]), .A2(n3743), .B1(rs1_val_gpr_w[27]), 
        .B2(n3376), .ZN(n3748) );
  NOR2_X1 U3958 ( .A1(rs2_val_gpr_w[24]), .A2(n3744), .ZN(n3745) );
  AOI22_X1 U3959 ( .A1(rs1_val_gpr_w[24]), .A2(n3745), .B1(rs1_val_gpr_w[25]), 
        .B2(n3384), .ZN(n3747) );
  AOI221_X1 U3960 ( .B1(n3759), .B2(n3748), .C1(n3747), .C2(n3748), .A(n3761), 
        .ZN(n3751) );
  OAI21_X1 U3961 ( .B1(rs1_val_gpr_w[31]), .B2(n3298), .A(rs1_val_gpr_w[30]), 
        .ZN(n3749) );
  OAI22_X1 U3962 ( .A1(rs2_val_gpr_w[30]), .A2(n3749), .B1(rs2_val_gpr_w[31]), 
        .B2(n3345), .ZN(n3750) );
  AOI211_X1 U3963 ( .C1(n3760), .C2(n3752), .A(n3751), .B(n3750), .ZN(n3753)
         );
  OAI221_X1 U3964 ( .B1(n3756), .B2(n3755), .C1(n3756), .C2(n3754), .A(n3753), 
        .ZN(u_branch_N127) );
  INV_X1 U3965 ( .A(n3684), .ZN(n3759) );
  INV_X1 U3966 ( .A(n3702), .ZN(n3757) );
  INV_X1 U3967 ( .A(n3724), .ZN(n3758) );
  INV_X1 U3968 ( .A(n3740), .ZN(n3760) );
  INV_X1 U3969 ( .A(n3746), .ZN(n3761) );
  XNOR2_X1 U3970 ( .A(rs1_val_gpr_w[31]), .B(mem_i_inst_i[31]), .ZN(n3762) );
  XNOR2_X1 U3971 ( .A(n3762), .B(add_x_67_n2), .ZN(mem_addr_w[31]) );
  NAND2_X1 U3972 ( .A1(n6581), .A2(n6577), .ZN(n6466) );
  AOI21_X1 U3973 ( .B1(u_branch_N120), .B2(n6741), .A(n6448), .ZN(n6454) );
  BUF_X1 U3974 ( .A(n5811), .Z(n4782) );
  NAND2_X1 U3975 ( .A1(n3520), .A2(mem_i_inst_i[15]), .ZN(n4942) );
  BUF_X1 U3976 ( .A(n7227), .Z(n4830) );
  BUF_X1 U3977 ( .A(n7251), .Z(n4831) );
  NOR3_X1 U3978 ( .A1(n7641), .A2(n7640), .A3(n7639), .ZN(n7642) );
  AOI211_X1 U3979 ( .C1(alu_b_q[28]), .C2(n7763), .A(n7762), .B(n7761), .ZN(
        n7764) );
  AOI22_X1 U3980 ( .A1(n7630), .A2(n7629), .B1(n3792), .B2(n3841), .ZN(n7655)
         );
  AOI21_X1 U3981 ( .B1(n7593), .B2(n7592), .A(n7591), .ZN(n7630) );
  AOI22_X1 U3982 ( .A1(n3766), .A2(n3839), .B1(n7575), .B2(n7574), .ZN(n7593)
         );
  AOI221_X1 U3983 ( .B1(n3775), .B2(n7293), .C1(n3813), .C2(n7293), .A(n7292), 
        .ZN(n7303) );
  AOI222_X1 U3984 ( .A1(alu_a_q[10]), .A2(alu_b_q[10]), .B1(alu_a_q[10]), .B2(
        n7252), .C1(alu_b_q[10]), .C2(n7252), .ZN(n7293) );
  OAI22_X1 U3985 ( .A1(n7117), .A2(n7116), .B1(n3809), .B2(n3780), .ZN(n7140)
         );
  AOI22_X1 U3986 ( .A1(alu_b_q[3]), .A2(alu_a_q[3]), .B1(n7095), .B2(n7094), 
        .ZN(n7116) );
  OAI22_X1 U3987 ( .A1(n7074), .A2(n7073), .B1(n3763), .B2(n3803), .ZN(n7094)
         );
  INV_X1 U3988 ( .A(n7054), .ZN(n7074) );
  NOR2_X1 U3989 ( .A1(n7731), .A2(n7930), .ZN(n7767) );
  NOR2_X1 U3990 ( .A1(n7718), .A2(n7889), .ZN(n7731) );
  AOI21_X1 U3991 ( .B1(alu_b_q[25]), .B2(n3829), .A(n7685), .ZN(n7718) );
  NAND2_X1 U3992 ( .A1(n7628), .A2(n7923), .ZN(n7645) );
  AOI22_X1 U3993 ( .A1(n7915), .A2(n7555), .B1(n3791), .B2(alu_b_q[20]), .ZN(
        n7576) );
  NAND2_X1 U3994 ( .A1(n7910), .A2(n7483), .ZN(n7509) );
  NAND2_X1 U3995 ( .A1(n7459), .A2(n7460), .ZN(n7483) );
  INV_X1 U3996 ( .A(n7289), .ZN(n7291) );
  NAND2_X1 U3997 ( .A1(n7253), .A2(n7899), .ZN(n7289) );
  OAI22_X1 U3998 ( .A1(alu_b_q[6]), .A2(n3773), .B1(n7163), .B2(n7162), .ZN(
        n7185) );
  AOI22_X1 U3999 ( .A1(alu_a_q[5]), .A2(n3812), .B1(n7139), .B2(n7138), .ZN(
        n7162) );
  OAI221_X1 U4000 ( .B1(n7119), .B2(alu_b_q[4]), .C1(n7119), .C2(n3780), .A(
        n7118), .ZN(n7138) );
  NAND2_X1 U4001 ( .A1(alu_b_q[0]), .A2(n3808), .ZN(n7068) );
  BUF_X1 U4002 ( .A(n7184), .Z(n4829) );
  BUF_X1 U4003 ( .A(n7161), .Z(n4828) );
  NOR2_X1 U4004 ( .A1(n7441), .A2(n7440), .ZN(n7442) );
  AOI211_X1 U4005 ( .C1(n7699), .C2(n7588), .A(n7587), .B(n7586), .ZN(n7589)
         );
  AOI211_X1 U4006 ( .C1(n3352), .C2(n7670), .A(n7669), .B(n7668), .ZN(n7671)
         );
  AOI22_X1 U4007 ( .A1(alu_a_q[26]), .A2(alu_b_q[26]), .B1(n7715), .B2(n7714), 
        .ZN(n7733) );
  OAI21_X1 U4008 ( .B1(alu_a_q[5]), .B2(alu_b_q[5]), .A(n7140), .ZN(n7141) );
  OAI22_X1 U4009 ( .A1(alu_b_q[1]), .A2(alu_a_q[1]), .B1(n7049), .B2(n7870), 
        .ZN(n7073) );
  INV_X1 U4010 ( .A(n7122), .ZN(n7146) );
  INV_X1 U4011 ( .A(n7883), .ZN(n7125) );
  OAI21_X1 U4012 ( .B1(n7767), .B2(n7888), .A(n7766), .ZN(n7813) );
  INV_X1 U4013 ( .A(n6786), .ZN(mem_i_rd_o) );
  OR2_X1 U4014 ( .A1(rst_i), .A2(n4821), .ZN(n3796) );
  INV_X1 U4015 ( .A(n6726), .ZN(n_1_net_) );
  BUF_X1 U4016 ( .A(n5811), .Z(n4779) );
  OAI22_X1 U4017 ( .A1(n6676), .A2(n6675), .B1(n6674), .B2(n6673), .ZN(
        mem_misaligned_w) );
  NOR2_X1 U4018 ( .A1(n4944), .A2(mem_i_inst_i[16]), .ZN(n6385) );
  INV_X1 U4019 ( .A(mem_i_inst_i[13]), .ZN(n6684) );
  INV_X1 U4020 ( .A(mem_i_inst_i[6]), .ZN(n6754) );
  INV_X1 U4021 ( .A(mem_i_inst_i[31]), .ZN(n4910) );
  BUF_X1 U4022 ( .A(n7007), .Z(n4824) );
  INV_X1 U4023 ( .A(n6678), .ZN(n6862) );
  AOI211_X1 U4024 ( .C1(n7519), .C2(n7518), .A(n7517), .B(n7516), .ZN(n7520)
         );
  AOI211_X1 U4025 ( .C1(n7739), .C2(n7544), .A(n7543), .B(n7542), .ZN(n7545)
         );
  NOR4_X1 U4026 ( .A1(n7613), .A2(n7612), .A3(n7611), .A4(n7610), .ZN(n7614)
         );
  INV_X1 U4027 ( .A(n7831), .ZN(n7699) );
  INV_X1 U4028 ( .A(n7342), .ZN(n7735) );
  BUF_X1 U4029 ( .A(n7975), .Z(n4889) );
  BUF_X1 U4030 ( .A(n7976), .Z(n4891) );
  BUF_X1 U4031 ( .A(n7980), .Z(n4899) );
  BUF_X1 U4032 ( .A(n7979), .Z(n4897) );
  BUF_X1 U4033 ( .A(n7978), .Z(n4895) );
  BUF_X1 U4034 ( .A(n7977), .Z(n4893) );
  INV_X1 U4035 ( .A(n7399), .ZN(n7425) );
  BUF_X1 U4036 ( .A(n7981), .Z(n4901) );
  BUF_X1 U4037 ( .A(n7971), .Z(n4881) );
  BUF_X1 U4038 ( .A(n7968), .Z(n4875) );
  BUF_X1 U4039 ( .A(n7967), .Z(n4873) );
  BUF_X1 U4040 ( .A(n7984), .Z(n4907) );
  BUF_X1 U4041 ( .A(n7983), .Z(n4905) );
  BUF_X1 U4042 ( .A(n7974), .Z(n4887) );
  BUF_X1 U4043 ( .A(n7985), .Z(n4909) );
  BUF_X1 U4044 ( .A(n7962), .Z(n4863) );
  BUF_X1 U4045 ( .A(n7961), .Z(n4861) );
  BUF_X1 U4046 ( .A(n7973), .Z(n4885) );
  BUF_X1 U4047 ( .A(n7972), .Z(n4883) );
  BUF_X1 U4048 ( .A(n7958), .Z(n4855) );
  BUF_X1 U4049 ( .A(n7963), .Z(n4865) );
  BUF_X1 U4050 ( .A(n7956), .Z(n4851) );
  BUF_X1 U4051 ( .A(n7982), .Z(n4903) );
  BUF_X1 U4052 ( .A(n7954), .Z(n4847) );
  BUF_X1 U4053 ( .A(n7970), .Z(n4879) );
  BUF_X1 U4054 ( .A(n7955), .Z(n4849) );
  BUF_X1 U4055 ( .A(n7957), .Z(n4853) );
  BUF_X1 U4056 ( .A(n7965), .Z(n4869) );
  BUF_X1 U4057 ( .A(n7964), .Z(n4867) );
  BUF_X1 U4058 ( .A(n7966), .Z(n4871) );
  BUF_X1 U4059 ( .A(n7969), .Z(n4877) );
  BUF_X1 U4060 ( .A(n7959), .Z(n4857) );
  INV_X1 U4061 ( .A(n7734), .ZN(n7872) );
  AOI21_X1 U4062 ( .B1(n7818), .B2(n7817), .A(n7816), .ZN(n7853) );
  AOI22_X1 U4063 ( .A1(n7733), .A2(n7732), .B1(n3784), .B2(n3843), .ZN(n7769)
         );
  INV_X1 U4064 ( .A(n7101), .ZN(n7082) );
  INV_X1 U4065 ( .A(n7414), .ZN(n7427) );
  INV_X1 U4066 ( .A(n7865), .ZN(n7835) );
  INV_X1 U4067 ( .A(n7282), .ZN(n7424) );
  NOR2_X1 U4068 ( .A1(n7929), .A2(n7813), .ZN(n7829) );
  BUF_X1 U4069 ( .A(n7960), .Z(n4859) );
  AOI21_X1 U4070 ( .B1(n4819), .B2(n3297), .A(n6468), .ZN(n6559) );
  NAND2_X1 U4071 ( .A1(n6467), .A2(n6462), .ZN(n6577) );
  BUF_X1 U4072 ( .A(n6383), .Z(n4796) );
  BUF_X1 U4073 ( .A(n3799), .Z(n4777) );
  BUF_X1 U4074 ( .A(n3769), .Z(n4768) );
  INV_X1 U4075 ( .A(mem_i_inst_i[19]), .ZN(n6619) );
  INV_X1 U4076 ( .A(mem_i_inst_i[18]), .ZN(n6615) );
  OR4_X1 U4077 ( .A1(n6750), .A2(n6844), .A3(n6791), .A4(n6776), .ZN(n6788) );
  INV_X1 U4078 ( .A(mem_i_inst_i[12]), .ZN(n6685) );
  INV_X1 U4079 ( .A(mem_i_inst_i[4]), .ZN(n6755) );
  NOR2_X1 U4080 ( .A1(mem_i_inst_i[2]), .A2(mem_i_inst_i[3]), .ZN(n6756) );
  BUF_X1 U4081 ( .A(n7008), .Z(n4825) );
  BUF_X1 U4082 ( .A(n7006), .Z(n4823) );
  INV_X1 U4083 ( .A(n6838), .ZN(n6840) );
  NOR3_X1 U4084 ( .A1(n7250), .A2(n7249), .A3(n7248), .ZN(n7251) );
  AOI211_X1 U4085 ( .C1(n7364), .C2(n7363), .A(n7362), .B(n7361), .ZN(n7365)
         );
  AOI211_X1 U4086 ( .C1(n7336), .C2(n7331), .A(n7330), .B(n7329), .ZN(n7332)
         );
  NOR4_X1 U4087 ( .A1(n7566), .A2(n7565), .A3(n7564), .A4(n7563), .ZN(n7567)
         );
  INV_X1 U4088 ( .A(n7385), .ZN(n7874) );
  INV_X1 U4089 ( .A(n7389), .ZN(n7885) );
  NOR2_X1 U4090 ( .A1(n7046), .A2(n7041), .ZN(n7980) );
  NOR2_X1 U4091 ( .A1(n7046), .A2(n7040), .ZN(n7979) );
  NOR2_X1 U4092 ( .A1(n7046), .A2(n7039), .ZN(n7978) );
  INV_X1 U4093 ( .A(n7620), .ZN(n7808) );
  INV_X1 U4094 ( .A(n7707), .ZN(n7866) );
  INV_X1 U4095 ( .A(n7708), .ZN(n7801) );
  INV_X1 U4096 ( .A(n7833), .ZN(n7797) );
  INV_X1 U4097 ( .A(n7709), .ZN(n7796) );
  NOR2_X1 U4098 ( .A1(n7046), .A2(n7042), .ZN(n7981) );
  NOR2_X1 U4099 ( .A1(n7037), .A2(n7040), .ZN(n7971) );
  NOR2_X1 U4100 ( .A1(n7046), .A2(n7045), .ZN(n7984) );
  NOR2_X1 U4101 ( .A1(n7046), .A2(n7044), .ZN(n7983) );
  NOR2_X1 U4102 ( .A1(n7037), .A2(n7043), .ZN(n7974) );
  NOR2_X1 U4103 ( .A1(n7046), .A2(n7047), .ZN(n7985) );
  NOR2_X1 U4104 ( .A1(n7037), .A2(n7042), .ZN(n7973) );
  NOR2_X1 U4105 ( .A1(n7037), .A2(n7041), .ZN(n7972) );
  NOR2_X1 U4106 ( .A1(n7046), .A2(n7043), .ZN(n7982) );
  NAND2_X1 U4107 ( .A1(n7038), .A2(n3868), .ZN(n7046) );
  NOR2_X1 U4108 ( .A1(n7037), .A2(n7039), .ZN(n7970) );
  INV_X1 U4109 ( .A(n7660), .ZN(n7856) );
  AND2_X1 U4110 ( .A1(alu_a_q[14]), .A2(alu_b_q[14]), .ZN(n7369) );
  NOR2_X1 U4111 ( .A1(n3835), .A2(n7941), .ZN(n7887) );
  NAND2_X1 U4112 ( .A1(n3807), .A2(n3774), .ZN(n7774) );
  NOR2_X1 U4113 ( .A1(n6874), .A2(exception_w), .ZN(n6845) );
  INV_X1 U4114 ( .A(n6750), .ZN(n6743) );
  INV_X1 U4115 ( .A(n6461), .ZN(n6467) );
  BUF_X1 U4116 ( .A(n5811), .Z(n4778) );
  NAND2_X1 U4117 ( .A1(n6472), .A2(n6587), .ZN(n6551) );
  INV_X1 U4118 ( .A(rst_i), .ZN(n6877) );
  NAND4_X1 U4119 ( .A1(n6756), .A2(mem_i_inst_i[5]), .A3(n6755), .A4(n6754), 
        .ZN(n7990) );
  OR2_X1 U4120 ( .A1(mem_i_inst_i[23]), .A2(mem_i_inst_i[24]), .ZN(n3800) );
  INV_X1 U4121 ( .A(mem_i_inst_i[14]), .ZN(n6821) );
  NOR3_X1 U4122 ( .A1(mem_i_inst_i[30]), .A2(n6824), .A3(n6749), .ZN(n6750) );
  INV_X1 U4123 ( .A(mem_i_inst_i[3]), .ZN(n6686) );
  INV_X1 U4124 ( .A(mem_i_inst_i[26]), .ZN(n6827) );
  INV_X1 U4125 ( .A(mem_i_inst_i[27]), .ZN(n6830) );
  INV_X1 U4126 ( .A(mem_i_inst_i[25]), .ZN(n6824) );
  AND2_X1 U4127 ( .A1(n159), .A2(n6959), .ZN(n7005) );
  INV_X1 U4128 ( .A(n6925), .ZN(n6951) );
  INV_X1 U4129 ( .A(n6924), .ZN(n6952) );
  INV_X1 U4130 ( .A(n6918), .ZN(n4826) );
  NAND2_X1 U4131 ( .A1(n6773), .A2(n6772), .ZN(n6918) );
  AOI211_X1 U4132 ( .C1(n7183), .C2(n7186), .A(n7182), .B(n7181), .ZN(n7184)
         );
  AOI221_X1 U4133 ( .B1(n7835), .B2(n7160), .C1(n7159), .C2(n7160), .A(n7158), 
        .ZN(n7161) );
  INV_X1 U4134 ( .A(n6793), .ZN(n6813) );
  AOI211_X1 U4135 ( .C1(n7242), .C2(n7226), .A(n7225), .B(n7224), .ZN(n7227)
         );
  AOI211_X1 U4136 ( .C1(n7292), .C2(n7274), .A(n7273), .B(n7272), .ZN(n7275)
         );
  AOI211_X1 U4137 ( .C1(n7425), .C2(n7738), .A(n7300), .B(n7299), .ZN(n7301)
         );
  NOR4_X1 U4138 ( .A1(n7403), .A2(n7402), .A3(n7401), .A4(n7400), .ZN(n7404)
         );
  NOR4_X1 U4139 ( .A1(n7470), .A2(n7469), .A3(n7468), .A4(n7467), .ZN(n7471)
         );
  INV_X1 U4140 ( .A(n6866), .ZN(n6677) );
  NOR4_X1 U4141 ( .A1(n7493), .A2(n7492), .A3(n7491), .A4(n7490), .ZN(n7494)
         );
  AND4_X1 U4142 ( .A1(n6684), .A2(n6685), .A3(n6870), .A4(n6846), .ZN(n6858)
         );
  NOR4_X1 U4143 ( .A1(n7793), .A2(n7792), .A3(n7791), .A4(n7790), .ZN(n7794)
         );
  AND4_X1 U4144 ( .A1(n7525), .A2(n7524), .A3(n7523), .A4(n7522), .ZN(n7750)
         );
  INV_X2 U4145 ( .A(n4889), .ZN(n4888) );
  NOR2_X1 U4146 ( .A1(n7037), .A2(n7044), .ZN(n7975) );
  INV_X2 U4147 ( .A(n4891), .ZN(n4890) );
  NOR2_X1 U4148 ( .A1(n7037), .A2(n7045), .ZN(n7976) );
  INV_X2 U4149 ( .A(n4899), .ZN(n4898) );
  INV_X2 U4150 ( .A(n4897), .ZN(n4896) );
  INV_X2 U4151 ( .A(n4895), .ZN(n4894) );
  INV_X2 U4152 ( .A(n4893), .ZN(n4892) );
  NOR2_X1 U4153 ( .A1(n7037), .A2(n7047), .ZN(n7977) );
  NAND2_X1 U4154 ( .A1(n3830), .A2(n7856), .ZN(n7788) );
  NAND2_X1 U4155 ( .A1(n7414), .A2(n7425), .ZN(n7707) );
  NAND2_X1 U4156 ( .A1(n7846), .A2(n3809), .ZN(n7399) );
  INV_X2 U4157 ( .A(n4901), .ZN(n4900) );
  INV_X2 U4158 ( .A(n4881), .ZN(n4880) );
  INV_X2 U4159 ( .A(n4875), .ZN(n4874) );
  NOR2_X1 U4160 ( .A1(n7035), .A2(n7045), .ZN(n7968) );
  INV_X2 U4161 ( .A(n4873), .ZN(n4872) );
  NOR2_X1 U4162 ( .A1(n7035), .A2(n7044), .ZN(n7967) );
  INV_X2 U4163 ( .A(n4907), .ZN(n4906) );
  INV_X2 U4164 ( .A(n4905), .ZN(n4904) );
  INV_X2 U4165 ( .A(n4887), .ZN(n4886) );
  INV_X2 U4166 ( .A(n4909), .ZN(n4908) );
  INV_X2 U4167 ( .A(n4863), .ZN(n4862) );
  NOR2_X1 U4168 ( .A1(n7035), .A2(n7039), .ZN(n7962) );
  INV_X2 U4169 ( .A(n4861), .ZN(n4860) );
  NOR2_X1 U4170 ( .A1(n7034), .A2(n7047), .ZN(n7961) );
  INV_X2 U4171 ( .A(n4885), .ZN(n4884) );
  INV_X2 U4172 ( .A(n4883), .ZN(n4882) );
  INV_X2 U4173 ( .A(n4855), .ZN(n4854) );
  NOR2_X1 U4174 ( .A1(n7034), .A2(n7043), .ZN(n7958) );
  INV_X2 U4175 ( .A(n4865), .ZN(n4864) );
  NOR2_X1 U4176 ( .A1(n7035), .A2(n7040), .ZN(n7963) );
  INV_X2 U4177 ( .A(n4851), .ZN(n4850) );
  NOR2_X1 U4178 ( .A1(n7034), .A2(n7041), .ZN(n7956) );
  INV_X2 U4179 ( .A(n4903), .ZN(n4902) );
  INV_X2 U4180 ( .A(n4847), .ZN(n4846) );
  NOR2_X1 U4181 ( .A1(n7034), .A2(n7039), .ZN(n7954) );
  INV_X2 U4182 ( .A(n4879), .ZN(n4878) );
  NAND2_X1 U4183 ( .A1(n144), .A2(n7038), .ZN(n7037) );
  NOR2_X1 U4184 ( .A1(n143), .A2(n7036), .ZN(n7038) );
  INV_X2 U4185 ( .A(n4849), .ZN(n4848) );
  NOR2_X1 U4186 ( .A1(n7034), .A2(n7040), .ZN(n7955) );
  INV_X2 U4187 ( .A(n4853), .ZN(n4852) );
  NOR2_X1 U4188 ( .A1(n7034), .A2(n7042), .ZN(n7957) );
  INV_X2 U4189 ( .A(n4869), .ZN(n4868) );
  NOR2_X1 U4190 ( .A1(n7035), .A2(n7042), .ZN(n7965) );
  INV_X2 U4191 ( .A(n4867), .ZN(n4866) );
  NOR2_X1 U4192 ( .A1(n7035), .A2(n7041), .ZN(n7964) );
  INV_X2 U4193 ( .A(n4871), .ZN(n4870) );
  NOR2_X1 U4194 ( .A1(n7035), .A2(n7043), .ZN(n7966) );
  INV_X2 U4195 ( .A(n4877), .ZN(n4876) );
  NOR2_X1 U4196 ( .A1(n7035), .A2(n7047), .ZN(n7969) );
  NAND4_X1 U4197 ( .A1(n143), .A2(mem_i_rd_o), .A3(rd_wr_en_q), .A4(n3868), 
        .ZN(n7035) );
  INV_X2 U4198 ( .A(n4857), .ZN(n4856) );
  NOR2_X1 U4199 ( .A1(n7034), .A2(n7044), .ZN(n7959) );
  INV_X2 U4200 ( .A(n4859), .ZN(n4858) );
  NAND2_X1 U4201 ( .A1(n157), .A2(n7624), .ZN(n7734) );
  INV_X1 U4202 ( .A(n7417), .ZN(n7313) );
  NAND2_X1 U4203 ( .A1(n7887), .A2(n3809), .ZN(n7831) );
  NAND4_X1 U4204 ( .A1(n7864), .A2(n7660), .A3(n7941), .A4(n7025), .ZN(n7867)
         );
  NOR2_X1 U4205 ( .A1(n7430), .A2(n7429), .ZN(n7833) );
  NAND2_X1 U4206 ( .A1(alu_b_q[4]), .A2(n7887), .ZN(n7430) );
  NAND2_X1 U4207 ( .A1(n3830), .A2(n7624), .ZN(n7865) );
  NOR4_X1 U4208 ( .A1(n157), .A2(n3765), .A3(n3788), .A4(n3835), .ZN(n7846) );
  NOR2_X1 U4209 ( .A1(n3772), .A2(alu_b_q[2]), .ZN(n7417) );
  NAND2_X1 U4210 ( .A1(alu_b_q[1]), .A2(alu_b_q[0]), .ZN(n7122) );
  NAND2_X1 U4211 ( .A1(n3774), .A2(alu_b_q[1]), .ZN(n7883) );
  NOR2_X2 U4212 ( .A1(n3774), .A2(alu_b_q[1]), .ZN(n7101) );
  NAND3_X1 U4213 ( .A1(n3788), .A2(n157), .A3(n154), .ZN(n7864) );
  NOR2_X1 U4214 ( .A1(n7034), .A2(n7045), .ZN(n7960) );
  NAND4_X1 U4215 ( .A1(n144), .A2(n143), .A3(mem_i_rd_o), .A4(rd_wr_en_q), 
        .ZN(n7034) );
  NAND2_X1 U4216 ( .A1(n57), .A2(state_q_0_), .ZN(n6786) );
  NAND2_X1 U4217 ( .A1(n6683), .A2(mem_i_valid_i), .ZN(n6726) );
  AND2_X1 U4218 ( .A1(n6682), .A2(n6750), .ZN(inst_div_w) );
  INV_X1 U4219 ( .A(n6493), .ZN(n6554) );
  NOR2_X1 U4220 ( .A1(n6472), .A2(n6471), .ZN(n6589) );
  AND2_X1 U4221 ( .A1(mem_i_inst_i[14]), .A2(mem_i_inst_i[13]), .ZN(n6680) );
  BUF_X1 U4222 ( .A(n5805), .Z(n4754) );
  INV_X1 U4223 ( .A(n3800), .ZN(n4816) );
  INV_X1 U4224 ( .A(mem_i_inst_i[24]), .ZN(n6573) );
  INV_X1 U4225 ( .A(mem_i_inst_i[23]), .ZN(n6576) );
  INV_X1 U4226 ( .A(n6468), .ZN(n6587) );
  INV_X1 U4227 ( .A(n6874), .ZN(n6870) );
  NAND2_X1 U4228 ( .A1(mem_i_valid_i), .A2(n6877), .ZN(n6874) );
  INV_X1 U4229 ( .A(n6404), .ZN(n4817) );
  INV_X1 U4230 ( .A(mem_i_inst_i[8]), .ZN(n7988) );
  INV_X1 U4231 ( .A(n6835), .ZN(n6841) );
  INV_X1 U4232 ( .A(n6880), .ZN(n6637) );
  NAND2_X1 U4233 ( .A1(n6814), .A2(n6813), .ZN(n6880) );
  NOR3_X1 U4234 ( .A1(rst_i), .A2(n6878), .A3(n6876), .ZN(n7006) );
  AOI211_X1 U4235 ( .C1(alu_b_q[2]), .C2(n7067), .A(n7066), .B(n7065), .ZN(
        n5090) );
  AOI211_X1 U4236 ( .C1(n7033), .C2(n7887), .A(n7031), .B(n7032), .ZN(n5033)
         );
  NAND2_X1 U4237 ( .A1(n6792), .A2(n4824), .ZN(n6838) );
  NOR2_X1 U4238 ( .A1(n6791), .A2(n6793), .ZN(n7007) );
  AOI211_X1 U4239 ( .C1(alu_a_q[3]), .C2(n7802), .A(n7092), .B(n7091), .ZN(
        n7093) );
  AOI21_X1 U4240 ( .B1(n7136), .B2(n7135), .A(n7134), .ZN(n7137) );
  NAND2_X1 U4241 ( .A1(n6870), .A2(n6772), .ZN(n6793) );
  AND2_X1 U4242 ( .A1(n7914), .A2(n7530), .ZN(n7519) );
  INV_X1 U4243 ( .A(n7851), .ZN(n7739) );
  NAND3_X1 U4244 ( .A1(n147), .A2(n145), .A3(n146), .ZN(n7039) );
  NAND2_X1 U4245 ( .A1(mem_i_rd_o), .A2(rd_wr_en_q), .ZN(n7036) );
  NAND3_X1 U4246 ( .A1(n145), .A2(n146), .A3(n3798), .ZN(n7040) );
  NAND3_X1 U4247 ( .A1(n145), .A2(n3798), .A3(n3865), .ZN(n7042) );
  NAND3_X1 U4248 ( .A1(n145), .A2(n147), .A3(n3865), .ZN(n7041) );
  NAND3_X1 U4249 ( .A1(n147), .A2(n146), .A3(n3767), .ZN(n7043) );
  NAND3_X1 U4250 ( .A1(n3798), .A2(n3767), .A3(n3865), .ZN(n7047) );
  NAND3_X1 U4251 ( .A1(n146), .A2(n3798), .A3(n3767), .ZN(n7044) );
  NAND2_X1 U4252 ( .A1(alu_b_q[4]), .A2(n7846), .ZN(n7851) );
  NAND2_X1 U4253 ( .A1(n3772), .A2(alu_b_q[2]), .ZN(n7282) );
  NOR2_X1 U4254 ( .A1(n3772), .A2(n3763), .ZN(n7418) );
  NAND3_X1 U4255 ( .A1(n147), .A2(n3767), .A3(n3865), .ZN(n7045) );
  INV_X1 U4256 ( .A(n6680), .ZN(n6744) );
  NOR2_X1 U4257 ( .A1(rst_i), .A2(mem_i_valid_i), .ZN(n6773) );
  BUF_X1 U4258 ( .A(n6383), .Z(n4793) );
  BUF_X1 U4259 ( .A(n6383), .Z(n4794) );
  BUF_X1 U4260 ( .A(n6383), .Z(n4792) );
  BUF_X1 U4261 ( .A(n5811), .Z(n4784) );
  BUF_X1 U4262 ( .A(n3799), .Z(n4769) );
  BUF_X1 U4263 ( .A(n3769), .Z(n4761) );
  BUF_X1 U4264 ( .A(n3799), .Z(n4770) );
  BUF_X1 U4265 ( .A(n5811), .Z(n4785) );
  BUF_X1 U4266 ( .A(n3769), .Z(n4762) );
  BUF_X1 U4267 ( .A(n5810), .Z(n4760) );
  BUF_X1 U4268 ( .A(n6383), .Z(n4795) );
  NAND4_X1 U4269 ( .A1(n6362), .A2(n6361), .A3(n6360), .A4(n6359), .ZN(
        rs1_val_gpr_w[29]) );
  BUF_X1 U4270 ( .A(n6383), .Z(n4797) );
  INV_X1 U4271 ( .A(mem_i_inst_i[7]), .ZN(n7986) );
  NOR2_X1 U4272 ( .A1(mem_i_inst_i[19]), .A2(mem_i_inst_i[18]), .ZN(n6397) );
  NOR2_X2 U4273 ( .A1(n4910), .A2(n6811), .ZN(n6835) );
  NOR2_X2 U4274 ( .A1(n6853), .A2(n6855), .ZN(n6863) );
  NAND2_X1 U4275 ( .A1(n155), .A2(n3765), .ZN(n7941) );
  AOI211_X1 U4276 ( .C1(n7117), .C2(n7114), .A(n7113), .B(n7112), .ZN(n7115)
         );
  NOR2_X1 U4277 ( .A1(n6573), .A2(mem_i_inst_i[23]), .ZN(n5804) );
  NOR2_X1 U4278 ( .A1(n6576), .A2(mem_i_inst_i[24]), .ZN(n5808) );
  NOR2_X1 U4279 ( .A1(state_q_0_), .A2(n3837), .ZN(n6760) );
  OAI22_X1 U4280 ( .A1(n6673), .A2(n6874), .B1(n161), .B2(n6875), .ZN(n2812)
         );
  OAI22_X1 U4281 ( .A1(n6676), .A2(n6874), .B1(n160), .B2(n6875), .ZN(n2813)
         );
  INV_X1 U4282 ( .A(n6773), .ZN(n6875) );
  AOI21_X1 U4283 ( .B1(n6839), .B2(csr_data_w[2]), .A(n6409), .ZN(n6796) );
  OAI22_X1 U4284 ( .A1(n6838), .A2(n3309), .B1(n6811), .B2(n6410), .ZN(n6409)
         );
  OAI21_X1 U4285 ( .B1(n5090), .B2(n4890), .A(n5060), .ZN(n2724) );
  NAND2_X1 U4286 ( .A1(n4890), .A2(reg_file[290]), .ZN(n5060) );
  OAI21_X1 U4287 ( .B1(n5033), .B2(n4886), .A(n5004), .ZN(n2758) );
  NAND2_X1 U4288 ( .A1(n4886), .A2(reg_file[353]), .ZN(n5004) );
  OAI21_X1 U4289 ( .B1(n5033), .B2(n4890), .A(n5003), .ZN(n2756) );
  NAND2_X1 U4290 ( .A1(n4890), .A2(reg_file[289]), .ZN(n5003) );
  OAI21_X1 U4291 ( .B1(n5090), .B2(n4886), .A(n5061), .ZN(n2726) );
  NAND2_X1 U4292 ( .A1(n4886), .A2(reg_file[354]), .ZN(n5061) );
  OAI21_X1 U4293 ( .B1(n5090), .B2(n4878), .A(n5059), .ZN(n2730) );
  NAND2_X1 U4294 ( .A1(n4878), .A2(reg_file[482]), .ZN(n5059) );
  OAI21_X1 U4295 ( .B1(n5033), .B2(n4878), .A(n5002), .ZN(n2762) );
  NAND2_X1 U4296 ( .A1(n4878), .A2(reg_file[481]), .ZN(n5002) );
  OAI21_X1 U4297 ( .B1(n5090), .B2(n4880), .A(n5058), .ZN(n2729) );
  NAND2_X1 U4298 ( .A1(n4880), .A2(reg_file[450]), .ZN(n5058) );
  OAI21_X1 U4299 ( .B1(n5033), .B2(n4880), .A(n5001), .ZN(n2761) );
  NAND2_X1 U4300 ( .A1(n4880), .A2(reg_file[449]), .ZN(n5001) );
  OAI21_X1 U4301 ( .B1(n7093), .B2(n4868), .A(n5145), .ZN(n2703) );
  NAND2_X1 U4302 ( .A1(n4868), .A2(reg_file[643]), .ZN(n5145) );
  OAI21_X1 U4303 ( .B1(n7093), .B2(n4870), .A(n5142), .ZN(n2702) );
  NAND2_X1 U4304 ( .A1(n4870), .A2(reg_file[611]), .ZN(n5142) );
  OAI21_X1 U4305 ( .B1(n7093), .B2(n4866), .A(n5146), .ZN(n2704) );
  NAND2_X1 U4306 ( .A1(n4866), .A2(reg_file[675]), .ZN(n5146) );
  AOI22_X1 U4307 ( .A1(n4825), .A2(mem_i_pc_o[28]), .B1(n7007), .B2(
        rs1_val_gpr_w[28]), .ZN(n6997) );
  AOI22_X1 U4308 ( .A1(n4825), .A2(mem_i_pc_o[31]), .B1(n7007), .B2(
        rs1_val_gpr_w[31]), .ZN(n7010) );
  AOI22_X1 U4309 ( .A1(n4825), .A2(mem_i_pc_o[30]), .B1(n7007), .B2(
        rs1_val_gpr_w[30]), .ZN(n7003) );
  AOI22_X1 U4310 ( .A1(n4825), .A2(mem_i_pc_o[26]), .B1(n7007), .B2(
        rs1_val_gpr_w[26]), .ZN(n6991) );
  AOI22_X1 U4311 ( .A1(n4825), .A2(mem_i_pc_o[27]), .B1(n7007), .B2(
        rs1_val_gpr_w[27]), .ZN(n6994) );
  AOI22_X1 U4312 ( .A1(n4825), .A2(mem_i_pc_o[29]), .B1(n7007), .B2(
        rs1_val_gpr_w[29]), .ZN(n7000) );
  OAI21_X1 U4313 ( .B1(n3372), .B2(n4848), .A(n5195), .ZN(n2681) );
  NAND2_X1 U4314 ( .A1(n4848), .A2(reg_file[964]), .ZN(n5195) );
  OAI21_X1 U4315 ( .B1(n3372), .B2(n4846), .A(n5196), .ZN(n2682) );
  NAND2_X1 U4316 ( .A1(n4846), .A2(reg_file[996]), .ZN(n5196) );
  OAI21_X1 U4317 ( .B1(n3372), .B2(n4866), .A(n5186), .ZN(n2672) );
  NAND2_X1 U4318 ( .A1(n4866), .A2(reg_file[676]), .ZN(n5186) );
  OAI21_X1 U4319 ( .B1(n3372), .B2(n4872), .A(n5184), .ZN(n2669) );
  NAND2_X1 U4320 ( .A1(n4872), .A2(reg_file[580]), .ZN(n5184) );
  OAI21_X1 U4321 ( .B1(n3372), .B2(n4874), .A(n5181), .ZN(n2668) );
  NAND2_X1 U4322 ( .A1(n4874), .A2(reg_file[548]), .ZN(n5181) );
  OAI21_X1 U4323 ( .B1(n3372), .B2(n4896), .A(n5171), .ZN(n2657) );
  NAND2_X1 U4324 ( .A1(n4896), .A2(reg_file[196]), .ZN(n5171) );
  OAI21_X1 U4325 ( .B1(n3372), .B2(n4876), .A(n5183), .ZN(n2667) );
  NAND2_X1 U4326 ( .A1(n4876), .A2(reg_file[516]), .ZN(n5183) );
  OAI21_X1 U4327 ( .B1(n3372), .B2(n4908), .A(n5175), .ZN(n2651) );
  NAND2_X1 U4328 ( .A1(n4908), .A2(reg_file[4]), .ZN(n5175) );
  OAI21_X1 U4329 ( .B1(n3372), .B2(n4906), .A(n5173), .ZN(n2652) );
  NAND2_X1 U4330 ( .A1(n4906), .A2(reg_file[36]), .ZN(n5173) );
  OAI21_X1 U4331 ( .B1(n3372), .B2(n4904), .A(n5176), .ZN(n2653) );
  NAND2_X1 U4332 ( .A1(n4904), .A2(reg_file[68]), .ZN(n5176) );
  OAI21_X1 U4333 ( .B1(n3372), .B2(n4902), .A(n5174), .ZN(n2654) );
  NAND2_X1 U4334 ( .A1(n4902), .A2(reg_file[100]), .ZN(n5174) );
  OAI21_X1 U4335 ( .B1(n3372), .B2(n4900), .A(n5177), .ZN(n2655) );
  NAND2_X1 U4336 ( .A1(n4900), .A2(reg_file[132]), .ZN(n5177) );
  OAI21_X1 U4337 ( .B1(n3372), .B2(n4898), .A(n5178), .ZN(n2656) );
  NAND2_X1 U4338 ( .A1(n4898), .A2(reg_file[164]), .ZN(n5178) );
  OAI21_X1 U4339 ( .B1(n3372), .B2(n4868), .A(n5185), .ZN(n2671) );
  NAND2_X1 U4340 ( .A1(n4868), .A2(reg_file[644]), .ZN(n5185) );
  OAI21_X1 U4341 ( .B1(n3372), .B2(n4870), .A(n5182), .ZN(n2670) );
  NAND2_X1 U4342 ( .A1(n4870), .A2(reg_file[612]), .ZN(n5182) );
  OAI21_X1 U4343 ( .B1(n3372), .B2(n4856), .A(n5200), .ZN(n2677) );
  NAND2_X1 U4344 ( .A1(n4856), .A2(reg_file[836]), .ZN(n5200) );
  OAI21_X1 U4345 ( .B1(n3372), .B2(n4860), .A(n5199), .ZN(n2675) );
  NAND2_X1 U4346 ( .A1(n4860), .A2(reg_file[772]), .ZN(n5199) );
  OAI21_X1 U4347 ( .B1(n3372), .B2(n4864), .A(n5179), .ZN(n2673) );
  NAND2_X1 U4348 ( .A1(n4864), .A2(reg_file[708]), .ZN(n5179) );
  OAI21_X1 U4349 ( .B1(n3372), .B2(n4854), .A(n5198), .ZN(n2678) );
  NAND2_X1 U4350 ( .A1(n4854), .A2(reg_file[868]), .ZN(n5198) );
  OAI21_X1 U4351 ( .B1(n3372), .B2(n4890), .A(n5189), .ZN(n2660) );
  NAND2_X1 U4352 ( .A1(n4890), .A2(reg_file[292]), .ZN(n5189) );
  OAI21_X1 U4353 ( .B1(n3372), .B2(n4852), .A(n5201), .ZN(n2679) );
  NAND2_X1 U4354 ( .A1(n4852), .A2(reg_file[900]), .ZN(n5201) );
  OAI21_X1 U4355 ( .B1(n3372), .B2(n4884), .A(n5193), .ZN(n2663) );
  NAND2_X1 U4356 ( .A1(n4884), .A2(reg_file[388]), .ZN(n5193) );
  OAI21_X1 U4357 ( .B1(n3372), .B2(n4850), .A(n5202), .ZN(n2680) );
  NAND2_X1 U4358 ( .A1(n4850), .A2(reg_file[932]), .ZN(n5202) );
  OAI21_X1 U4359 ( .B1(n3372), .B2(n4858), .A(n5197), .ZN(n2676) );
  NAND2_X1 U4360 ( .A1(n4858), .A2(reg_file[804]), .ZN(n5197) );
  OAI21_X1 U4361 ( .B1(n3372), .B2(n4880), .A(n5187), .ZN(n2665) );
  NAND2_X1 U4362 ( .A1(n4880), .A2(reg_file[452]), .ZN(n5187) );
  OAI21_X1 U4363 ( .B1(n3372), .B2(n4878), .A(n5188), .ZN(n2666) );
  NAND2_X1 U4364 ( .A1(n4878), .A2(reg_file[484]), .ZN(n5188) );
  OAI21_X1 U4365 ( .B1(n3372), .B2(n4886), .A(n5190), .ZN(n2662) );
  NAND2_X1 U4366 ( .A1(n4886), .A2(reg_file[356]), .ZN(n5190) );
  OAI21_X1 U4367 ( .B1(n3372), .B2(n4888), .A(n5192), .ZN(n2661) );
  NAND2_X1 U4368 ( .A1(n4888), .A2(reg_file[324]), .ZN(n5192) );
  OAI21_X1 U4369 ( .B1(n3372), .B2(n4892), .A(n5191), .ZN(n2659) );
  NAND2_X1 U4370 ( .A1(n4892), .A2(reg_file[260]), .ZN(n5191) );
  OAI21_X1 U4371 ( .B1(n3372), .B2(n4862), .A(n5180), .ZN(n2674) );
  NAND2_X1 U4372 ( .A1(n4862), .A2(reg_file[740]), .ZN(n5180) );
  OAI21_X1 U4373 ( .B1(n3372), .B2(n4894), .A(n5172), .ZN(n2658) );
  NAND2_X1 U4374 ( .A1(n4894), .A2(reg_file[228]), .ZN(n5172) );
  OAI21_X1 U4375 ( .B1(n3372), .B2(n4882), .A(n5194), .ZN(n2664) );
  NAND2_X1 U4376 ( .A1(n4882), .A2(reg_file[420]), .ZN(n5194) );
  OAI21_X1 U4377 ( .B1(n3374), .B2(n4862), .A(n5083), .ZN(n2738) );
  NAND2_X1 U4378 ( .A1(n4862), .A2(reg_file[738]), .ZN(n5083) );
  OAI21_X1 U4379 ( .B1(n3374), .B2(n4884), .A(n5064), .ZN(n2727) );
  NAND2_X1 U4380 ( .A1(n4884), .A2(reg_file[386]), .ZN(n5064) );
  OAI21_X1 U4381 ( .B1(n3374), .B2(n4866), .A(n5089), .ZN(n2736) );
  NAND2_X1 U4382 ( .A1(n4866), .A2(reg_file[674]), .ZN(n5089) );
  OAI21_X1 U4383 ( .B1(n3374), .B2(n4876), .A(n5086), .ZN(n2731) );
  NAND2_X1 U4384 ( .A1(n4876), .A2(reg_file[514]), .ZN(n5086) );
  OAI21_X1 U4385 ( .B1(n3374), .B2(n4882), .A(n5065), .ZN(n2728) );
  NAND2_X1 U4386 ( .A1(n4882), .A2(reg_file[418]), .ZN(n5065) );
  OAI21_X1 U4387 ( .B1(n3374), .B2(n4872), .A(n5087), .ZN(n2733) );
  NAND2_X1 U4388 ( .A1(n4872), .A2(reg_file[578]), .ZN(n5087) );
  OAI21_X1 U4389 ( .B1(n3374), .B2(n4870), .A(n5085), .ZN(n2734) );
  NAND2_X1 U4390 ( .A1(n4870), .A2(reg_file[610]), .ZN(n5085) );
  OAI21_X1 U4391 ( .B1(n3374), .B2(n4874), .A(n5084), .ZN(n2732) );
  NAND2_X1 U4392 ( .A1(n4874), .A2(reg_file[546]), .ZN(n5084) );
  OAI21_X1 U4393 ( .B1(n3374), .B2(n4892), .A(n5062), .ZN(n2723) );
  NAND2_X1 U4394 ( .A1(n4892), .A2(reg_file[258]), .ZN(n5062) );
  OAI21_X1 U4395 ( .B1(n3374), .B2(n4868), .A(n5088), .ZN(n2735) );
  NAND2_X1 U4396 ( .A1(n4868), .A2(reg_file[642]), .ZN(n5088) );
  OAI21_X1 U4397 ( .B1(n3374), .B2(n4864), .A(n5082), .ZN(n2737) );
  NAND2_X1 U4398 ( .A1(n4864), .A2(reg_file[706]), .ZN(n5082) );
  OAI21_X1 U4399 ( .B1(n3375), .B2(n4850), .A(n5032), .ZN(n2776) );
  NAND2_X1 U4400 ( .A1(n4850), .A2(reg_file[929]), .ZN(n5032) );
  OAI21_X1 U4401 ( .B1(n3375), .B2(n4846), .A(n5026), .ZN(n2778) );
  NAND2_X1 U4402 ( .A1(n4846), .A2(reg_file[993]), .ZN(n5026) );
  OAI21_X1 U4403 ( .B1(n3375), .B2(n4852), .A(n5031), .ZN(n2775) );
  NAND2_X1 U4404 ( .A1(n4852), .A2(reg_file[897]), .ZN(n5031) );
  OAI21_X1 U4405 ( .B1(n3375), .B2(n4848), .A(n5025), .ZN(n2777) );
  NAND2_X1 U4406 ( .A1(n4848), .A2(reg_file[961]), .ZN(n5025) );
  OAI21_X1 U4407 ( .B1(n3375), .B2(n4882), .A(n5008), .ZN(n2760) );
  NAND2_X1 U4408 ( .A1(n4882), .A2(reg_file[417]), .ZN(n5008) );
  OAI21_X1 U4409 ( .B1(n3375), .B2(n4884), .A(n5007), .ZN(n2759) );
  NAND2_X1 U4410 ( .A1(n4884), .A2(reg_file[385]), .ZN(n5007) );
  OAI21_X1 U4411 ( .B1(n3375), .B2(n4858), .A(n5027), .ZN(n2772) );
  NAND2_X1 U4412 ( .A1(n4858), .A2(reg_file[801]), .ZN(n5027) );
  OAI21_X1 U4413 ( .B1(n3375), .B2(n4856), .A(n5030), .ZN(n2773) );
  NAND2_X1 U4414 ( .A1(n4856), .A2(reg_file[833]), .ZN(n5030) );
  OAI21_X1 U4415 ( .B1(n3375), .B2(n4854), .A(n5028), .ZN(n2774) );
  NAND2_X1 U4416 ( .A1(n4854), .A2(reg_file[865]), .ZN(n5028) );
  OAI21_X1 U4417 ( .B1(n3375), .B2(n4892), .A(n5005), .ZN(n2755) );
  NAND2_X1 U4418 ( .A1(n4892), .A2(reg_file[257]), .ZN(n5005) );
  OAI21_X1 U4419 ( .B1(n3375), .B2(n4860), .A(n5029), .ZN(n2771) );
  NAND2_X1 U4420 ( .A1(n4860), .A2(reg_file[769]), .ZN(n5029) );
  OAI21_X1 U4421 ( .B1(n7137), .B2(n4854), .A(n5248), .ZN(n2646) );
  NAND2_X1 U4422 ( .A1(n4854), .A2(reg_file[869]), .ZN(n5248) );
  OAI21_X1 U4423 ( .B1(n7137), .B2(n4860), .A(n5249), .ZN(n2643) );
  NAND2_X1 U4424 ( .A1(n4860), .A2(reg_file[773]), .ZN(n5249) );
  OAI21_X1 U4425 ( .B1(n7137), .B2(n4858), .A(n5247), .ZN(n2644) );
  NAND2_X1 U4426 ( .A1(n4858), .A2(reg_file[805]), .ZN(n5247) );
  OAI21_X1 U4427 ( .B1(n7137), .B2(n4856), .A(n5250), .ZN(n2645) );
  NAND2_X1 U4428 ( .A1(n4856), .A2(reg_file[837]), .ZN(n5250) );
  OAI21_X1 U4429 ( .B1(n7137), .B2(n4850), .A(n5252), .ZN(n2648) );
  NAND2_X1 U4430 ( .A1(n4850), .A2(reg_file[933]), .ZN(n5252) );
  OAI21_X1 U4431 ( .B1(n7137), .B2(n4852), .A(n5251), .ZN(n2647) );
  NAND2_X1 U4432 ( .A1(n4852), .A2(reg_file[901]), .ZN(n5251) );
  OAI21_X1 U4433 ( .B1(n6918), .B2(n3803), .A(n6898), .ZN(n6594) );
  OAI21_X1 U4434 ( .B1(n6918), .B2(n3779), .A(n6894), .ZN(n6598) );
  OAI211_X1 U4435 ( .C1(n3325), .C2(n6838), .A(n6665), .B(n6798), .ZN(n2870)
         );
  NAND2_X1 U4436 ( .A1(csr_data_w[4]), .A2(n6839), .ZN(n6665) );
  OAI211_X1 U4437 ( .C1(n3336), .C2(n6838), .A(n6639), .B(n6638), .ZN(n2850)
         );
  AOI211_X1 U4438 ( .C1(n6637), .C2(mem_i_inst_i[24]), .A(n6835), .B(n6636), 
        .ZN(n6638) );
  NOR2_X1 U4439 ( .A1(n3840), .A2(n6918), .ZN(n6636) );
  NAND2_X1 U4440 ( .A1(csr_data_w[24]), .A2(n6839), .ZN(n6639) );
  OAI211_X1 U4441 ( .C1(n3340), .C2(n6838), .A(n6614), .B(n6613), .ZN(n2857)
         );
  AOI211_X1 U4442 ( .C1(n4826), .C2(alu_b_q[17]), .A(n6835), .B(n6612), .ZN(
        n6613) );
  NOR2_X1 U4443 ( .A1(n6880), .A2(n3520), .ZN(n6612) );
  NAND2_X1 U4444 ( .A1(csr_data_w[17]), .A2(n6839), .ZN(n6614) );
  OAI211_X1 U4445 ( .C1(n3312), .C2(n6838), .A(n6629), .B(n6628), .ZN(n2853)
         );
  AOI211_X1 U4446 ( .C1(n6637), .C2(mem_i_inst_i[21]), .A(n6835), .B(n6627), 
        .ZN(n6628) );
  NOR2_X1 U4447 ( .A1(n3839), .A2(n6918), .ZN(n6627) );
  NAND2_X1 U4448 ( .A1(csr_data_w[21]), .A2(n6839), .ZN(n6629) );
  OAI211_X1 U4449 ( .C1(n3332), .C2(n6838), .A(n6622), .B(n6621), .ZN(n2855)
         );
  AOI211_X1 U4450 ( .C1(n4826), .C2(alu_b_q[19]), .A(n6835), .B(n6620), .ZN(
        n6621) );
  NOR2_X1 U4451 ( .A1(n6880), .A2(n6619), .ZN(n6620) );
  NAND2_X1 U4452 ( .A1(csr_data_w[19]), .A2(n6839), .ZN(n6622) );
  OAI211_X1 U4453 ( .C1(n3326), .C2(n6838), .A(n6626), .B(n6625), .ZN(n2854)
         );
  AOI211_X1 U4454 ( .C1(n4826), .C2(alu_b_q[20]), .A(n6835), .B(n6624), .ZN(
        n6625) );
  NOR2_X1 U4455 ( .A1(n6880), .A2(n6623), .ZN(n6624) );
  NAND2_X1 U4456 ( .A1(csr_data_w[20]), .A2(n6839), .ZN(n6626) );
  OAI211_X1 U4457 ( .C1(n3343), .C2(n6838), .A(n6632), .B(n6631), .ZN(n2852)
         );
  AOI211_X1 U4458 ( .C1(n6637), .C2(mem_i_inst_i[22]), .A(n6835), .B(n6630), 
        .ZN(n6631) );
  NOR2_X1 U4459 ( .A1(n3845), .A2(n6918), .ZN(n6630) );
  NAND2_X1 U4460 ( .A1(csr_data_w[22]), .A2(n6839), .ZN(n6632) );
  OAI211_X1 U4461 ( .C1(n3338), .C2(n6838), .A(n6611), .B(n6610), .ZN(n2858)
         );
  AOI211_X1 U4462 ( .C1(n4826), .C2(alu_b_q[16]), .A(n6835), .B(n6609), .ZN(
        n6610) );
  NOR2_X1 U4463 ( .A1(n6880), .A2(n6608), .ZN(n6609) );
  NAND2_X1 U4464 ( .A1(csr_data_w[16]), .A2(n6839), .ZN(n6611) );
  OAI211_X1 U4465 ( .C1(n3311), .C2(n6838), .A(n6607), .B(n6606), .ZN(n2859)
         );
  AOI211_X1 U4466 ( .C1(alu_b_q[15]), .C2(n4826), .A(n6835), .B(n6605), .ZN(
        n6606) );
  NOR2_X1 U4467 ( .A1(n6880), .A2(n6604), .ZN(n6605) );
  NAND2_X1 U4468 ( .A1(csr_data_w[15]), .A2(n6839), .ZN(n6607) );
  OAI211_X1 U4469 ( .C1(n3310), .C2(n6838), .A(n6635), .B(n6634), .ZN(n2851)
         );
  AOI211_X1 U4470 ( .C1(n6637), .C2(mem_i_inst_i[23]), .A(n6835), .B(n6633), 
        .ZN(n6634) );
  NOR2_X1 U4471 ( .A1(n3841), .A2(n6918), .ZN(n6633) );
  NAND2_X1 U4472 ( .A1(csr_data_w[23]), .A2(n6839), .ZN(n6635) );
  OAI211_X1 U4473 ( .C1(n3337), .C2(n6838), .A(n6618), .B(n6617), .ZN(n2856)
         );
  AOI211_X1 U4474 ( .C1(n4826), .C2(alu_b_q[18]), .A(n6835), .B(n6616), .ZN(
        n6617) );
  NOR2_X1 U4475 ( .A1(n6880), .A2(n6615), .ZN(n6616) );
  NAND2_X1 U4476 ( .A1(csr_data_w[18]), .A2(n6839), .ZN(n6618) );
  OAI211_X1 U4477 ( .C1(n3303), .C2(n6838), .A(n6664), .B(n6799), .ZN(n2869)
         );
  NAND2_X1 U4478 ( .A1(csr_data_w[5]), .A2(n6839), .ZN(n6664) );
  AOI211_X1 U4479 ( .C1(n4824), .C2(n3521), .A(n4970), .B(n6889), .ZN(n4971)
         );
  OAI21_X1 U4480 ( .B1(n6918), .B2(n3808), .A(n6890), .ZN(n4970) );
  AOI211_X1 U4481 ( .C1(n4824), .C2(n3524), .A(n6600), .B(n6901), .ZN(n6601)
         );
  OAI21_X1 U4482 ( .B1(n6918), .B2(n3804), .A(n6902), .ZN(n6600) );
  AOI211_X1 U4483 ( .C1(n4824), .C2(rs1_val_gpr_w[5]), .A(n6602), .B(n6909), 
        .ZN(n6603) );
  OAI21_X1 U4484 ( .B1(n6918), .B2(n3781), .A(n6910), .ZN(n6602) );
  AOI211_X1 U4485 ( .C1(n4824), .C2(rs1_val_gpr_w[4]), .A(n6596), .B(n6905), 
        .ZN(n6597) );
  OAI21_X1 U4486 ( .B1(n6918), .B2(n3780), .A(n6906), .ZN(n6596) );
  OAI21_X1 U4487 ( .B1(n3374), .B2(n4906), .A(n5076), .ZN(n2716) );
  NAND2_X1 U4488 ( .A1(n4906), .A2(reg_file[34]), .ZN(n5076) );
  OAI21_X1 U4489 ( .B1(n3374), .B2(n4902), .A(n5077), .ZN(n2718) );
  NAND2_X1 U4490 ( .A1(n4902), .A2(reg_file[98]), .ZN(n5077) );
  OAI21_X1 U4491 ( .B1(n3374), .B2(n4888), .A(n5063), .ZN(n2725) );
  NAND2_X1 U4492 ( .A1(n4888), .A2(reg_file[322]), .ZN(n5063) );
  OAI21_X1 U4493 ( .B1(n3374), .B2(n4896), .A(n5074), .ZN(n2721) );
  NAND2_X1 U4494 ( .A1(n4896), .A2(reg_file[194]), .ZN(n5074) );
  OAI21_X1 U4495 ( .B1(n3374), .B2(n4904), .A(n5079), .ZN(n2717) );
  NAND2_X1 U4496 ( .A1(n4904), .A2(reg_file[66]), .ZN(n5079) );
  OAI21_X1 U4497 ( .B1(n3374), .B2(n4908), .A(n5078), .ZN(n2715) );
  NAND2_X1 U4498 ( .A1(n4908), .A2(reg_file[2]), .ZN(n5078) );
  OAI21_X1 U4499 ( .B1(n3374), .B2(n4900), .A(n5080), .ZN(n2719) );
  NAND2_X1 U4500 ( .A1(n4900), .A2(reg_file[130]), .ZN(n5080) );
  OAI21_X1 U4501 ( .B1(n3374), .B2(n4894), .A(n5075), .ZN(n2722) );
  NAND2_X1 U4502 ( .A1(n4894), .A2(reg_file[226]), .ZN(n5075) );
  OAI21_X1 U4503 ( .B1(n3374), .B2(n4898), .A(n5081), .ZN(n2720) );
  NAND2_X1 U4504 ( .A1(n4898), .A2(reg_file[162]), .ZN(n5081) );
  OAI21_X1 U4505 ( .B1(n3374), .B2(n4858), .A(n5068), .ZN(n2740) );
  NAND2_X1 U4506 ( .A1(n4858), .A2(reg_file[802]), .ZN(n5068) );
  OAI21_X1 U4507 ( .B1(n3374), .B2(n4860), .A(n5070), .ZN(n2739) );
  NAND2_X1 U4508 ( .A1(n4860), .A2(reg_file[770]), .ZN(n5070) );
  OAI21_X1 U4509 ( .B1(n3374), .B2(n4846), .A(n5067), .ZN(n2746) );
  NAND2_X1 U4510 ( .A1(n4846), .A2(reg_file[994]), .ZN(n5067) );
  OAI21_X1 U4511 ( .B1(n3374), .B2(n4856), .A(n5071), .ZN(n2741) );
  NAND2_X1 U4512 ( .A1(n4856), .A2(reg_file[834]), .ZN(n5071) );
  OAI21_X1 U4513 ( .B1(n3374), .B2(n4854), .A(n5069), .ZN(n2742) );
  NAND2_X1 U4514 ( .A1(n4854), .A2(reg_file[866]), .ZN(n5069) );
  OAI21_X1 U4515 ( .B1(n3374), .B2(n4852), .A(n5072), .ZN(n2743) );
  NAND2_X1 U4516 ( .A1(n4852), .A2(reg_file[898]), .ZN(n5072) );
  OAI21_X1 U4517 ( .B1(n3374), .B2(n4850), .A(n5073), .ZN(n2744) );
  NAND2_X1 U4518 ( .A1(n4850), .A2(reg_file[930]), .ZN(n5073) );
  OAI21_X1 U4519 ( .B1(n3374), .B2(n4848), .A(n5066), .ZN(n2745) );
  NAND2_X1 U4520 ( .A1(n4848), .A2(reg_file[962]), .ZN(n5066) );
  OAI21_X1 U4521 ( .B1(n3375), .B2(n4900), .A(n5023), .ZN(n2751) );
  NAND2_X1 U4522 ( .A1(n4900), .A2(reg_file[129]), .ZN(n5023) );
  OAI21_X1 U4523 ( .B1(n3375), .B2(n4902), .A(n5020), .ZN(n2750) );
  NAND2_X1 U4524 ( .A1(n4902), .A2(reg_file[97]), .ZN(n5020) );
  OAI21_X1 U4525 ( .B1(n3375), .B2(n4888), .A(n5006), .ZN(n2757) );
  NAND2_X1 U4526 ( .A1(n4888), .A2(reg_file[321]), .ZN(n5006) );
  OAI21_X1 U4527 ( .B1(n3375), .B2(n4866), .A(n5016), .ZN(n2768) );
  NAND2_X1 U4528 ( .A1(n4866), .A2(reg_file[673]), .ZN(n5016) );
  OAI21_X1 U4529 ( .B1(n3375), .B2(n4894), .A(n5018), .ZN(n2754) );
  NAND2_X1 U4530 ( .A1(n4894), .A2(reg_file[225]), .ZN(n5018) );
  OAI21_X1 U4531 ( .B1(n3375), .B2(n4896), .A(n5017), .ZN(n2753) );
  NAND2_X1 U4532 ( .A1(n4896), .A2(reg_file[193]), .ZN(n5017) );
  OAI21_X1 U4533 ( .B1(n3375), .B2(n4898), .A(n5024), .ZN(n2752) );
  NAND2_X1 U4534 ( .A1(n4898), .A2(reg_file[161]), .ZN(n5024) );
  OAI21_X1 U4535 ( .B1(n3375), .B2(n4874), .A(n5011), .ZN(n2764) );
  NAND2_X1 U4536 ( .A1(n4874), .A2(reg_file[545]), .ZN(n5011) );
  OAI21_X1 U4537 ( .B1(n3375), .B2(n4876), .A(n5013), .ZN(n2763) );
  NAND2_X1 U4538 ( .A1(n4876), .A2(reg_file[513]), .ZN(n5013) );
  OAI21_X1 U4539 ( .B1(n3375), .B2(n4862), .A(n5010), .ZN(n2770) );
  NAND2_X1 U4540 ( .A1(n4862), .A2(reg_file[737]), .ZN(n5010) );
  OAI21_X1 U4541 ( .B1(n3375), .B2(n4864), .A(n5009), .ZN(n2769) );
  NAND2_X1 U4542 ( .A1(n4864), .A2(reg_file[705]), .ZN(n5009) );
  OAI21_X1 U4543 ( .B1(n3375), .B2(n4904), .A(n5022), .ZN(n2749) );
  NAND2_X1 U4544 ( .A1(n4904), .A2(reg_file[65]), .ZN(n5022) );
  OAI21_X1 U4545 ( .B1(n3375), .B2(n4868), .A(n5015), .ZN(n2767) );
  NAND2_X1 U4546 ( .A1(n4868), .A2(reg_file[641]), .ZN(n5015) );
  OAI21_X1 U4547 ( .B1(n3375), .B2(n4870), .A(n5012), .ZN(n2766) );
  NAND2_X1 U4548 ( .A1(n4870), .A2(reg_file[609]), .ZN(n5012) );
  OAI21_X1 U4549 ( .B1(n3375), .B2(n4872), .A(n5014), .ZN(n2765) );
  NAND2_X1 U4550 ( .A1(n4872), .A2(reg_file[577]), .ZN(n5014) );
  OAI21_X1 U4551 ( .B1(n3375), .B2(n4908), .A(n5021), .ZN(n2747) );
  NAND2_X1 U4552 ( .A1(n4908), .A2(reg_file[1]), .ZN(n5021) );
  OAI21_X1 U4553 ( .B1(n3375), .B2(n4906), .A(n5019), .ZN(n2748) );
  NAND2_X1 U4554 ( .A1(n4906), .A2(reg_file[33]), .ZN(n5019) );
  AOI21_X1 U4555 ( .B1(csr_data_w[3]), .B2(n6839), .A(n6666), .ZN(n6667) );
  OAI21_X1 U4556 ( .B1(n3299), .B2(n6838), .A(n6797), .ZN(n6666) );
  AOI21_X1 U4557 ( .B1(csr_data_w[1]), .B2(n6839), .A(n6668), .ZN(n6669) );
  OAI21_X1 U4558 ( .B1(n3302), .B2(n6838), .A(n6795), .ZN(n6668) );
  AOI21_X1 U4559 ( .B1(csr_data_w[0]), .B2(n6839), .A(n6670), .ZN(n6671) );
  OAI21_X1 U4560 ( .B1(n3328), .B2(n6838), .A(n6794), .ZN(n6670) );
  NOR2_X1 U4561 ( .A1(n6793), .A2(n6792), .ZN(n6808) );
  OAI21_X1 U4562 ( .B1(n3373), .B2(n4878), .A(n5116), .ZN(n2698) );
  NAND2_X1 U4563 ( .A1(n4878), .A2(reg_file[483]), .ZN(n5116) );
  OAI21_X1 U4564 ( .B1(n3373), .B2(n4880), .A(n5115), .ZN(n2697) );
  NAND2_X1 U4565 ( .A1(n4880), .A2(reg_file[451]), .ZN(n5115) );
  OAI21_X1 U4566 ( .B1(n3373), .B2(n4882), .A(n5122), .ZN(n2696) );
  NAND2_X1 U4567 ( .A1(n4882), .A2(reg_file[419]), .ZN(n5122) );
  OAI21_X1 U4568 ( .B1(n3373), .B2(n4846), .A(n5124), .ZN(n2714) );
  NAND2_X1 U4569 ( .A1(n4846), .A2(reg_file[995]), .ZN(n5124) );
  OAI21_X1 U4570 ( .B1(n3373), .B2(n4858), .A(n5125), .ZN(n2708) );
  NAND2_X1 U4571 ( .A1(n4858), .A2(reg_file[803]), .ZN(n5125) );
  OAI21_X1 U4572 ( .B1(n3373), .B2(n4888), .A(n5120), .ZN(n2693) );
  NAND2_X1 U4573 ( .A1(n4888), .A2(reg_file[323]), .ZN(n5120) );
  OAI21_X1 U4574 ( .B1(n3373), .B2(n4876), .A(n5143), .ZN(n2699) );
  NAND2_X1 U4575 ( .A1(n4876), .A2(reg_file[515]), .ZN(n5143) );
  OAI21_X1 U4576 ( .B1(n3373), .B2(n4854), .A(n5126), .ZN(n2710) );
  NAND2_X1 U4577 ( .A1(n4854), .A2(reg_file[867]), .ZN(n5126) );
  OAI21_X1 U4578 ( .B1(n3373), .B2(n4886), .A(n5118), .ZN(n2694) );
  NAND2_X1 U4579 ( .A1(n4886), .A2(reg_file[355]), .ZN(n5118) );
  OAI21_X1 U4580 ( .B1(n3373), .B2(n4884), .A(n5121), .ZN(n2695) );
  NAND2_X1 U4581 ( .A1(n4884), .A2(reg_file[387]), .ZN(n5121) );
  OAI21_X1 U4582 ( .B1(n3373), .B2(n4862), .A(n5140), .ZN(n2706) );
  NAND2_X1 U4583 ( .A1(n4862), .A2(reg_file[739]), .ZN(n5140) );
  OAI21_X1 U4584 ( .B1(n3373), .B2(n4892), .A(n5119), .ZN(n2691) );
  NAND2_X1 U4585 ( .A1(n4892), .A2(reg_file[259]), .ZN(n5119) );
  OAI21_X1 U4586 ( .B1(n3373), .B2(n4890), .A(n5117), .ZN(n2692) );
  NAND2_X1 U4587 ( .A1(n4890), .A2(reg_file[291]), .ZN(n5117) );
  OAI21_X1 U4588 ( .B1(n3373), .B2(n4848), .A(n5123), .ZN(n2713) );
  NAND2_X1 U4589 ( .A1(n4848), .A2(reg_file[963]), .ZN(n5123) );
  OAI21_X1 U4590 ( .B1(n3373), .B2(n4902), .A(n5134), .ZN(n2686) );
  NAND2_X1 U4591 ( .A1(n4902), .A2(reg_file[99]), .ZN(n5134) );
  OAI21_X1 U4592 ( .B1(n3373), .B2(n4856), .A(n5128), .ZN(n2709) );
  NAND2_X1 U4593 ( .A1(n4856), .A2(reg_file[835]), .ZN(n5128) );
  OAI21_X1 U4594 ( .B1(n3373), .B2(n4900), .A(n5137), .ZN(n2687) );
  NAND2_X1 U4595 ( .A1(n4900), .A2(reg_file[131]), .ZN(n5137) );
  OAI21_X1 U4596 ( .B1(n3373), .B2(n4908), .A(n5135), .ZN(n2683) );
  NAND2_X1 U4597 ( .A1(n4908), .A2(reg_file[3]), .ZN(n5135) );
  OAI21_X1 U4598 ( .B1(n3373), .B2(n4872), .A(n5144), .ZN(n2701) );
  NAND2_X1 U4599 ( .A1(n4872), .A2(reg_file[579]), .ZN(n5144) );
  OAI21_X1 U4600 ( .B1(n3373), .B2(n4874), .A(n5141), .ZN(n2700) );
  NAND2_X1 U4601 ( .A1(n4874), .A2(reg_file[547]), .ZN(n5141) );
  OAI21_X1 U4602 ( .B1(n3373), .B2(n4850), .A(n5130), .ZN(n2712) );
  NAND2_X1 U4603 ( .A1(n4850), .A2(reg_file[931]), .ZN(n5130) );
  OAI21_X1 U4604 ( .B1(n3373), .B2(n4860), .A(n5127), .ZN(n2707) );
  NAND2_X1 U4605 ( .A1(n4860), .A2(reg_file[771]), .ZN(n5127) );
  OAI21_X1 U4606 ( .B1(n3373), .B2(n4896), .A(n5131), .ZN(n2689) );
  NAND2_X1 U4607 ( .A1(n4896), .A2(reg_file[195]), .ZN(n5131) );
  OAI21_X1 U4608 ( .B1(n3373), .B2(n4852), .A(n5129), .ZN(n2711) );
  NAND2_X1 U4609 ( .A1(n4852), .A2(reg_file[899]), .ZN(n5129) );
  OAI21_X1 U4610 ( .B1(n3373), .B2(n4894), .A(n5132), .ZN(n2690) );
  NAND2_X1 U4611 ( .A1(n4894), .A2(reg_file[227]), .ZN(n5132) );
  OAI21_X1 U4612 ( .B1(n3373), .B2(n4898), .A(n5138), .ZN(n2688) );
  NAND2_X1 U4613 ( .A1(n4898), .A2(reg_file[163]), .ZN(n5138) );
  OAI21_X1 U4614 ( .B1(n3373), .B2(n4864), .A(n5139), .ZN(n2705) );
  NAND2_X1 U4615 ( .A1(n4864), .A2(reg_file[707]), .ZN(n5139) );
  OAI21_X1 U4616 ( .B1(n3373), .B2(n4904), .A(n5136), .ZN(n2685) );
  NAND2_X1 U4617 ( .A1(n4904), .A2(reg_file[67]), .ZN(n5136) );
  OAI21_X1 U4618 ( .B1(n3373), .B2(n4906), .A(n5133), .ZN(n2684) );
  NAND2_X1 U4619 ( .A1(n4906), .A2(reg_file[35]), .ZN(n5133) );
  OAI21_X1 U4620 ( .B1(n3371), .B2(n4878), .A(n5222), .ZN(n2634) );
  NAND2_X1 U4621 ( .A1(n4878), .A2(reg_file[485]), .ZN(n5222) );
  OAI21_X1 U4622 ( .B1(n3371), .B2(n4862), .A(n5230), .ZN(n2642) );
  NAND2_X1 U4623 ( .A1(n4862), .A2(reg_file[741]), .ZN(n5230) );
  OAI21_X1 U4624 ( .B1(n3371), .B2(n4848), .A(n5245), .ZN(n2649) );
  NAND2_X1 U4625 ( .A1(n4848), .A2(reg_file[965]), .ZN(n5245) );
  OAI21_X1 U4626 ( .B1(n3371), .B2(n4868), .A(n5235), .ZN(n2639) );
  NAND2_X1 U4627 ( .A1(n4868), .A2(reg_file[645]), .ZN(n5235) );
  OAI21_X1 U4628 ( .B1(n3371), .B2(n4904), .A(n5242), .ZN(n2621) );
  NAND2_X1 U4629 ( .A1(n4904), .A2(reg_file[69]), .ZN(n5242) );
  OAI21_X1 U4630 ( .B1(n3371), .B2(n4906), .A(n5239), .ZN(n2620) );
  NAND2_X1 U4631 ( .A1(n4906), .A2(reg_file[37]), .ZN(n5239) );
  OAI21_X1 U4632 ( .B1(n3371), .B2(n4866), .A(n5236), .ZN(n2640) );
  NAND2_X1 U4633 ( .A1(n4866), .A2(reg_file[677]), .ZN(n5236) );
  OAI21_X1 U4634 ( .B1(n3371), .B2(n4908), .A(n5241), .ZN(n2619) );
  NAND2_X1 U4635 ( .A1(n4908), .A2(reg_file[5]), .ZN(n5241) );
  OAI21_X1 U4636 ( .B1(n3371), .B2(n4896), .A(n5237), .ZN(n2625) );
  NAND2_X1 U4637 ( .A1(n4896), .A2(reg_file[197]), .ZN(n5237) );
  OAI21_X1 U4638 ( .B1(n3371), .B2(n4898), .A(n5244), .ZN(n2624) );
  NAND2_X1 U4639 ( .A1(n4898), .A2(reg_file[165]), .ZN(n5244) );
  OAI21_X1 U4640 ( .B1(n3371), .B2(n4900), .A(n5243), .ZN(n2623) );
  NAND2_X1 U4641 ( .A1(n4900), .A2(reg_file[133]), .ZN(n5243) );
  OAI21_X1 U4642 ( .B1(n3371), .B2(n4902), .A(n5240), .ZN(n2622) );
  NAND2_X1 U4643 ( .A1(n4902), .A2(reg_file[101]), .ZN(n5240) );
  OAI21_X1 U4644 ( .B1(n3371), .B2(n4884), .A(n5227), .ZN(n2631) );
  NAND2_X1 U4645 ( .A1(n4884), .A2(reg_file[389]), .ZN(n5227) );
  OAI21_X1 U4646 ( .B1(n3371), .B2(n4886), .A(n5224), .ZN(n2630) );
  NAND2_X1 U4647 ( .A1(n4886), .A2(reg_file[357]), .ZN(n5224) );
  OAI21_X1 U4648 ( .B1(n3371), .B2(n4888), .A(n5226), .ZN(n2629) );
  NAND2_X1 U4649 ( .A1(n4888), .A2(reg_file[325]), .ZN(n5226) );
  OAI21_X1 U4650 ( .B1(n3371), .B2(n4890), .A(n5223), .ZN(n2628) );
  NAND2_X1 U4651 ( .A1(n4890), .A2(reg_file[293]), .ZN(n5223) );
  OAI21_X1 U4652 ( .B1(n3371), .B2(n4892), .A(n5225), .ZN(n2627) );
  NAND2_X1 U4653 ( .A1(n4892), .A2(reg_file[261]), .ZN(n5225) );
  OAI21_X1 U4654 ( .B1(n3371), .B2(n4894), .A(n5238), .ZN(n2626) );
  NAND2_X1 U4655 ( .A1(n4894), .A2(reg_file[229]), .ZN(n5238) );
  OAI21_X1 U4656 ( .B1(n3371), .B2(n4864), .A(n5229), .ZN(n2641) );
  NAND2_X1 U4657 ( .A1(n4864), .A2(reg_file[709]), .ZN(n5229) );
  OAI21_X1 U4658 ( .B1(n3371), .B2(n4882), .A(n5228), .ZN(n2632) );
  NAND2_X1 U4659 ( .A1(n4882), .A2(reg_file[421]), .ZN(n5228) );
  OAI21_X1 U4660 ( .B1(n3371), .B2(n4846), .A(n5246), .ZN(n2650) );
  NAND2_X1 U4661 ( .A1(n4846), .A2(reg_file[997]), .ZN(n5246) );
  OAI21_X1 U4662 ( .B1(n3371), .B2(n4874), .A(n5231), .ZN(n2636) );
  NAND2_X1 U4663 ( .A1(n4874), .A2(reg_file[549]), .ZN(n5231) );
  OAI21_X1 U4664 ( .B1(n3371), .B2(n4876), .A(n5233), .ZN(n2635) );
  NAND2_X1 U4665 ( .A1(n4876), .A2(reg_file[517]), .ZN(n5233) );
  OAI21_X1 U4666 ( .B1(n3371), .B2(n4870), .A(n5232), .ZN(n2638) );
  NAND2_X1 U4667 ( .A1(n4870), .A2(reg_file[613]), .ZN(n5232) );
  OAI21_X1 U4668 ( .B1(n3371), .B2(n4880), .A(n5221), .ZN(n2633) );
  NAND2_X1 U4669 ( .A1(n4880), .A2(reg_file[453]), .ZN(n5221) );
  OAI21_X1 U4670 ( .B1(n3371), .B2(n4872), .A(n5234), .ZN(n2637) );
  NAND2_X1 U4671 ( .A1(n4872), .A2(reg_file[581]), .ZN(n5234) );
  NOR2_X1 U4672 ( .A1(n7342), .A2(n7226), .ZN(n4752) );
  AOI22_X1 U4673 ( .A1(mem_addr_w[7]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[7]), .ZN(n1437) );
  AOI22_X1 U4674 ( .A1(mem_addr_w[10]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[10]), .ZN(n1440) );
  AOI22_X1 U4675 ( .A1(mem_addr_w[9]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[9]), .ZN(n1439) );
  AOI22_X1 U4676 ( .A1(mem_addr_w[2]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[2]), .ZN(n1432) );
  AOI22_X1 U4677 ( .A1(mem_addr_w[3]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[3]), .ZN(n1433) );
  AOI22_X1 U4678 ( .A1(mem_addr_w[4]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[4]), .ZN(n1434) );
  AOI22_X1 U4679 ( .A1(mem_addr_w[5]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[5]), .ZN(n1435) );
  AOI22_X1 U4680 ( .A1(mem_addr_w[6]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[6]), .ZN(n1436) );
  AOI22_X1 U4681 ( .A1(mem_addr_w[8]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[8]), .ZN(n1438) );
  AOI22_X1 U4682 ( .A1(mem_addr_w[11]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[11]), .ZN(n1441) );
  OAI21_X1 U4683 ( .B1(n6862), .B2(n3328), .A(n6646), .ZN(n2827) );
  AOI22_X1 U4684 ( .A1(rs2_val_gpr_w[16]), .A2(n6863), .B1(n4822), .B2(
        mem_d_data_wr_o[16]), .ZN(n6646) );
  OAI21_X1 U4685 ( .B1(n6862), .B2(n3309), .A(n6648), .ZN(n2829) );
  AOI22_X1 U4686 ( .A1(rs2_val_gpr_w[18]), .A2(n6863), .B1(n4822), .B2(
        mem_d_data_wr_o[18]), .ZN(n6648) );
  OAI21_X1 U4687 ( .B1(n6862), .B2(n3325), .A(n6650), .ZN(n2831) );
  AOI22_X1 U4688 ( .A1(rs2_val_gpr_w[20]), .A2(n6863), .B1(n4822), .B2(
        mem_d_data_wr_o[20]), .ZN(n6650) );
  OAI21_X1 U4689 ( .B1(n6862), .B2(n3302), .A(n6647), .ZN(n2828) );
  AOI22_X1 U4690 ( .A1(rs2_val_gpr_w[17]), .A2(n6863), .B1(n4822), .B2(
        mem_d_data_wr_o[17]), .ZN(n6647) );
  OAI21_X1 U4691 ( .B1(n6862), .B2(n3299), .A(n6649), .ZN(n2830) );
  AOI22_X1 U4692 ( .A1(rs2_val_gpr_w[19]), .A2(n6863), .B1(n4822), .B2(
        mem_d_data_wr_o[19]), .ZN(n6649) );
  OAI21_X1 U4693 ( .B1(n6862), .B2(n3303), .A(n6651), .ZN(n2832) );
  AOI22_X1 U4694 ( .A1(rs2_val_gpr_w[21]), .A2(n6863), .B1(n4822), .B2(
        mem_d_data_wr_o[21]), .ZN(n6651) );
  OAI21_X1 U4695 ( .B1(n6865), .B2(n3325), .A(n6644), .ZN(n2823) );
  AOI22_X1 U4696 ( .A1(n6677), .A2(rs2_val_gpr_w[12]), .B1(n4822), .B2(
        mem_d_data_wr_o[12]), .ZN(n6644) );
  OAI21_X1 U4697 ( .B1(n6865), .B2(n3299), .A(n6643), .ZN(n2822) );
  AOI22_X1 U4698 ( .A1(n6677), .A2(rs2_val_gpr_w[11]), .B1(n4822), .B2(
        mem_d_data_wr_o[11]), .ZN(n6643) );
  OAI21_X1 U4699 ( .B1(n6865), .B2(n3303), .A(n6645), .ZN(n2824) );
  AOI22_X1 U4700 ( .A1(n6677), .A2(rs2_val_gpr_w[13]), .B1(n4822), .B2(
        mem_d_data_wr_o[13]), .ZN(n6645) );
  OAI21_X1 U4701 ( .B1(n6865), .B2(n3328), .A(n6640), .ZN(n2819) );
  AOI22_X1 U4702 ( .A1(n6677), .A2(rs2_val_gpr_w[8]), .B1(n4822), .B2(
        mem_d_data_wr_o[8]), .ZN(n6640) );
  OAI21_X1 U4703 ( .B1(n6865), .B2(n3302), .A(n6641), .ZN(n2820) );
  AOI22_X1 U4704 ( .A1(n6677), .A2(rs2_val_gpr_w[9]), .B1(n4822), .B2(
        mem_d_data_wr_o[9]), .ZN(n6641) );
  OAI21_X1 U4705 ( .B1(n6865), .B2(n3309), .A(n6642), .ZN(n2821) );
  AOI22_X1 U4706 ( .A1(n6677), .A2(rs2_val_gpr_w[10]), .B1(n4822), .B2(
        mem_d_data_wr_o[10]), .ZN(n6642) );
  NAND3_X1 U4707 ( .A1(n6858), .A2(mem_addr_w[0]), .A3(n6676), .ZN(n6865) );
  AOI22_X1 U4708 ( .A1(n6868), .A2(rs2_val_gpr_w[3]), .B1(n4822), .B2(
        mem_d_data_wr_o[3]), .ZN(n1383) );
  AOI22_X1 U4709 ( .A1(n6868), .A2(rs2_val_gpr_w[2]), .B1(n4822), .B2(
        mem_d_data_wr_o[2]), .ZN(n1382) );
  AOI22_X1 U4710 ( .A1(n6868), .A2(rs2_val_gpr_w[5]), .B1(n4822), .B2(
        mem_d_data_wr_o[5]), .ZN(n1385) );
  AOI22_X1 U4711 ( .A1(n6868), .A2(rs2_val_gpr_w[4]), .B1(n4822), .B2(
        mem_d_data_wr_o[4]), .ZN(n1384) );
  NAND2_X1 U4712 ( .A1(n6414), .A2(n6866), .ZN(n6868) );
  NAND3_X1 U4713 ( .A1(n6858), .A2(n6676), .A3(n6673), .ZN(n6414) );
  AOI22_X1 U4714 ( .A1(mem_addr_w[12]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[12]), .ZN(n1442) );
  AOI22_X1 U4715 ( .A1(mem_addr_w[13]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[13]), .ZN(n1443) );
  OAI211_X1 U4716 ( .C1(n6860), .C2(n3309), .A(n6657), .B(n6656), .ZN(n2837)
         );
  NAND2_X1 U4717 ( .A1(rs2_val_gpr_w[26]), .A2(n6863), .ZN(n6656) );
  AOI22_X1 U4718 ( .A1(rs2_val_gpr_w[10]), .A2(n6859), .B1(n4822), .B2(
        mem_d_data_wr_o[26]), .ZN(n6657) );
  OAI211_X1 U4719 ( .C1(n6860), .C2(n3328), .A(n6653), .B(n6652), .ZN(n2835)
         );
  NAND2_X1 U4720 ( .A1(rs2_val_gpr_w[24]), .A2(n6863), .ZN(n6652) );
  AOI22_X1 U4721 ( .A1(rs2_val_gpr_w[8]), .A2(n6859), .B1(n4822), .B2(
        mem_d_data_wr_o[24]), .ZN(n6653) );
  OAI211_X1 U4722 ( .C1(n6860), .C2(n3302), .A(n6655), .B(n6654), .ZN(n2836)
         );
  NAND2_X1 U4723 ( .A1(rs2_val_gpr_w[25]), .A2(n6863), .ZN(n6654) );
  AOI22_X1 U4724 ( .A1(rs2_val_gpr_w[9]), .A2(n6859), .B1(n4822), .B2(
        mem_d_data_wr_o[25]), .ZN(n6655) );
  OAI211_X1 U4725 ( .C1(n6860), .C2(n3303), .A(n6663), .B(n6662), .ZN(n2840)
         );
  NAND2_X1 U4726 ( .A1(rs2_val_gpr_w[29]), .A2(n6863), .ZN(n6662) );
  AOI22_X1 U4727 ( .A1(rs2_val_gpr_w[13]), .A2(n6859), .B1(n4822), .B2(
        mem_d_data_wr_o[29]), .ZN(n6663) );
  OAI211_X1 U4728 ( .C1(n6860), .C2(n3325), .A(n6661), .B(n6660), .ZN(n2839)
         );
  NAND2_X1 U4729 ( .A1(rs2_val_gpr_w[28]), .A2(n6863), .ZN(n6660) );
  AOI22_X1 U4730 ( .A1(rs2_val_gpr_w[12]), .A2(n6859), .B1(n4822), .B2(
        mem_d_data_wr_o[28]), .ZN(n6661) );
  OAI211_X1 U4731 ( .C1(n6860), .C2(n3299), .A(n6659), .B(n6658), .ZN(n2838)
         );
  NAND2_X1 U4732 ( .A1(rs2_val_gpr_w[27]), .A2(n6863), .ZN(n6658) );
  AOI22_X1 U4733 ( .A1(rs2_val_gpr_w[11]), .A2(n6859), .B1(n4822), .B2(
        mem_d_data_wr_o[27]), .ZN(n6659) );
  NOR2_X1 U4734 ( .A1(n6413), .A2(n6412), .ZN(n6678) );
  INV_X1 U4735 ( .A(n6846), .ZN(n6412) );
  NAND2_X1 U4736 ( .A1(mem_addr_w[1]), .A2(n6673), .ZN(n6413) );
  NAND3_X1 U4737 ( .A1(n6858), .A2(mem_addr_w[1]), .A3(mem_addr_w[0]), .ZN(
        n6860) );
  AOI22_X1 U4738 ( .A1(mem_addr_w[14]), .A2(n6845), .B1(n4822), .B2(
        mem_d_addr_o[14]), .ZN(n1444) );
  AOI22_X1 U4739 ( .A1(mem_addr_w[15]), .A2(n6845), .B1(n4822), .B2(
        mem_d_addr_o[15]), .ZN(n1445) );
  AOI22_X1 U4740 ( .A1(mem_addr_w[16]), .A2(n6845), .B1(n4822), .B2(
        mem_d_addr_o[16]), .ZN(n1446) );
  AOI22_X1 U4741 ( .A1(mem_addr_w[17]), .A2(n6845), .B1(n4822), .B2(
        mem_d_addr_o[17]), .ZN(n1447) );
  AOI22_X1 U4742 ( .A1(mem_addr_w[18]), .A2(n6845), .B1(n4822), .B2(
        mem_d_addr_o[18]), .ZN(n1448) );
  AOI22_X1 U4743 ( .A1(mem_addr_w[19]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[19]), .ZN(n1449) );
  OAI21_X1 U4744 ( .B1(n4973), .B2(n4874), .A(n4915), .ZN(n1772) );
  NAND2_X1 U4745 ( .A1(n4874), .A2(reg_file[544]), .ZN(n4915) );
  OAI21_X1 U4746 ( .B1(n4973), .B2(n4866), .A(n4911), .ZN(n1776) );
  NAND2_X1 U4747 ( .A1(n4866), .A2(reg_file[672]), .ZN(n4911) );
  OAI21_X1 U4748 ( .B1(n4973), .B2(n4870), .A(n4914), .ZN(n1774) );
  NAND2_X1 U4749 ( .A1(n4870), .A2(reg_file[608]), .ZN(n4914) );
  OAI21_X1 U4750 ( .B1(n4973), .B2(n4872), .A(n4913), .ZN(n1773) );
  NAND2_X1 U4751 ( .A1(n4872), .A2(reg_file[576]), .ZN(n4913) );
  OAI21_X1 U4752 ( .B1(n4973), .B2(n4864), .A(n4912), .ZN(n1777) );
  NAND2_X1 U4753 ( .A1(n4864), .A2(reg_file[704]), .ZN(n4912) );
  AOI22_X1 U4754 ( .A1(mem_addr_w[20]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[20]), .ZN(n1450) );
  OAI21_X1 U4755 ( .B1(n4973), .B2(n4848), .A(n4935), .ZN(n1785) );
  NAND2_X1 U4756 ( .A1(n4848), .A2(reg_file[960]), .ZN(n4935) );
  OAI21_X1 U4757 ( .B1(n4973), .B2(n4854), .A(n4937), .ZN(n1782) );
  NAND2_X1 U4758 ( .A1(n4854), .A2(reg_file[864]), .ZN(n4937) );
  OAI21_X1 U4759 ( .B1(n4973), .B2(n4868), .A(n4916), .ZN(n1775) );
  NAND2_X1 U4760 ( .A1(n4868), .A2(reg_file[640]), .ZN(n4916) );
  OAI21_X1 U4761 ( .B1(n4973), .B2(n4856), .A(n4936), .ZN(n1781) );
  NAND2_X1 U4762 ( .A1(n4856), .A2(reg_file[832]), .ZN(n4936) );
  OAI21_X1 U4763 ( .B1(n4973), .B2(n4846), .A(n4941), .ZN(n1786) );
  NAND2_X1 U4764 ( .A1(n4846), .A2(reg_file[992]), .ZN(n4941) );
  OAI21_X1 U4765 ( .B1(n4973), .B2(n4852), .A(n4939), .ZN(n1783) );
  NAND2_X1 U4766 ( .A1(n4852), .A2(reg_file[896]), .ZN(n4939) );
  OAI21_X1 U4767 ( .B1(n4973), .B2(n4860), .A(n4940), .ZN(n1779) );
  NAND2_X1 U4768 ( .A1(n4860), .A2(reg_file[768]), .ZN(n4940) );
  OAI21_X1 U4769 ( .B1(n4973), .B2(n4896), .A(n4972), .ZN(n1761) );
  NAND2_X1 U4770 ( .A1(n4896), .A2(reg_file[192]), .ZN(n4972) );
  OAI21_X1 U4771 ( .B1(n4973), .B2(n4862), .A(n4918), .ZN(n1778) );
  NAND2_X1 U4772 ( .A1(n4862), .A2(reg_file[736]), .ZN(n4918) );
  OAI21_X1 U4773 ( .B1(n4973), .B2(n4858), .A(n4938), .ZN(n1780) );
  NAND2_X1 U4774 ( .A1(n4858), .A2(reg_file[800]), .ZN(n4938) );
  OAI21_X1 U4775 ( .B1(n4753), .B2(n4904), .A(n4928), .ZN(n1757) );
  NAND2_X1 U4776 ( .A1(n4904), .A2(reg_file[64]), .ZN(n4928) );
  OAI21_X1 U4777 ( .B1(n4753), .B2(n4902), .A(n4929), .ZN(n1758) );
  NAND2_X1 U4778 ( .A1(n4902), .A2(reg_file[96]), .ZN(n4929) );
  OAI21_X1 U4779 ( .B1(n4753), .B2(n4900), .A(n4931), .ZN(n1759) );
  NAND2_X1 U4780 ( .A1(n4900), .A2(reg_file[128]), .ZN(n4931) );
  OAI21_X1 U4781 ( .B1(n4753), .B2(n4898), .A(n4927), .ZN(n1760) );
  NAND2_X1 U4782 ( .A1(n4898), .A2(reg_file[160]), .ZN(n4927) );
  OAI21_X1 U4783 ( .B1(n4753), .B2(n4894), .A(n4933), .ZN(n1762) );
  NAND2_X1 U4784 ( .A1(n4894), .A2(reg_file[224]), .ZN(n4933) );
  OAI21_X1 U4785 ( .B1(n4753), .B2(n4892), .A(n4925), .ZN(n1763) );
  NAND2_X1 U4786 ( .A1(n4892), .A2(reg_file[256]), .ZN(n4925) );
  OAI21_X1 U4787 ( .B1(n4753), .B2(n4890), .A(n4923), .ZN(n1764) );
  NAND2_X1 U4788 ( .A1(n4890), .A2(reg_file[288]), .ZN(n4923) );
  OAI21_X1 U4789 ( .B1(n4753), .B2(n4888), .A(n4921), .ZN(n1765) );
  NAND2_X1 U4790 ( .A1(n4888), .A2(reg_file[320]), .ZN(n4921) );
  OAI21_X1 U4791 ( .B1(n4753), .B2(n4886), .A(n4922), .ZN(n1766) );
  NAND2_X1 U4792 ( .A1(n4886), .A2(reg_file[352]), .ZN(n4922) );
  OAI21_X1 U4793 ( .B1(n4753), .B2(n4884), .A(n4924), .ZN(n1767) );
  NAND2_X1 U4794 ( .A1(n4884), .A2(reg_file[384]), .ZN(n4924) );
  OAI21_X1 U4795 ( .B1(n4753), .B2(n4882), .A(n4919), .ZN(n1768) );
  NAND2_X1 U4796 ( .A1(n4882), .A2(reg_file[416]), .ZN(n4919) );
  OAI21_X1 U4797 ( .B1(n4753), .B2(n4908), .A(n4932), .ZN(n1755) );
  NAND2_X1 U4798 ( .A1(n4908), .A2(reg_file[0]), .ZN(n4932) );
  OAI21_X1 U4799 ( .B1(n4753), .B2(n4880), .A(n4920), .ZN(n1769) );
  NAND2_X1 U4800 ( .A1(n4880), .A2(reg_file[448]), .ZN(n4920) );
  OAI21_X1 U4801 ( .B1(n4753), .B2(n4878), .A(n4926), .ZN(n1770) );
  NAND2_X1 U4802 ( .A1(n4878), .A2(reg_file[480]), .ZN(n4926) );
  OAI21_X1 U4803 ( .B1(n4753), .B2(n4876), .A(n4917), .ZN(n1771) );
  NAND2_X1 U4804 ( .A1(n4876), .A2(reg_file[512]), .ZN(n4917) );
  OAI21_X1 U4805 ( .B1(n4753), .B2(n4850), .A(n4934), .ZN(n1784) );
  NAND2_X1 U4806 ( .A1(n4850), .A2(reg_file[928]), .ZN(n4934) );
  OAI21_X1 U4807 ( .B1(n4753), .B2(n4906), .A(n4930), .ZN(n1756) );
  NAND2_X1 U4808 ( .A1(n4906), .A2(reg_file[32]), .ZN(n4930) );
  AOI22_X1 U4809 ( .A1(mem_addr_w[21]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[21]), .ZN(n1451) );
  OAI211_X1 U4810 ( .C1(n6593), .C2(n6592), .A(n6591), .B(n6590), .ZN(n2916)
         );
  AOI22_X1 U4811 ( .A1(n3319), .A2(csr_mepc_w[0]), .B1(n6588), .B2(
        mem_i_pc_o[0]), .ZN(n6590) );
  INV_X1 U4812 ( .A(reset_vector_i[0]), .ZN(n6592) );
  AOI22_X1 U4813 ( .A1(mem_addr_w[22]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[22]), .ZN(n1452) );
  AOI22_X1 U4814 ( .A1(mem_addr_w[23]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[23]), .ZN(n1453) );
  AOI22_X1 U4815 ( .A1(mem_addr_w[24]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[24]), .ZN(n1454) );
  INV_X1 U4816 ( .A(n6553), .ZN(n2912) );
  AOI21_X1 U4817 ( .B1(U4_RSOP_173_C3_DATA1_4), .B2(n6559), .A(n6552), .ZN(
        n6553) );
  OAI211_X1 U4818 ( .C1(reset_vector_i[4]), .C2(n6551), .A(n6550), .B(n6549), 
        .ZN(n6552) );
  AOI22_X1 U4819 ( .A1(n6588), .A2(mem_i_pc_o[4]), .B1(n6554), .B2(
        reset_vector_i[4]), .ZN(n6549) );
  NAND2_X1 U4820 ( .A1(n3319), .A2(csr_mepc_w[4]), .ZN(n6550) );
  AOI22_X1 U4821 ( .A1(mem_addr_w[25]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[25]), .ZN(n1455) );
  OAI211_X1 U4822 ( .C1(n6593), .C2(n6558), .A(n6557), .B(n6556), .ZN(n2913)
         );
  AOI22_X1 U4823 ( .A1(n3319), .A2(csr_mepc_w[3]), .B1(n6588), .B2(
        mem_i_pc_o[3]), .ZN(n6556) );
  NAND2_X1 U4824 ( .A1(U4_RSOP_173_C3_DATA1_3), .A2(n3363), .ZN(n6557) );
  INV_X1 U4825 ( .A(reset_vector_i[3]), .ZN(n6558) );
  NOR2_X1 U4826 ( .A1(n6555), .A2(n6554), .ZN(n6593) );
  AOI22_X1 U4827 ( .A1(mem_addr_w[26]), .A2(n6845), .B1(n4822), .B2(
        mem_d_addr_o[26]), .ZN(n1456) );
  AOI22_X1 U4828 ( .A1(mem_addr_w[27]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[27]), .ZN(n1457) );
  AOI22_X1 U4829 ( .A1(mem_addr_w[28]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[28]), .ZN(n1458) );
  INV_X1 U4830 ( .A(n6547), .ZN(n2908) );
  AOI21_X1 U4831 ( .B1(U4_RSOP_173_C3_DATA1_8), .B2(n6559), .A(n6546), .ZN(
        n6547) );
  OAI211_X1 U4832 ( .C1(n6761), .C2(n6551), .A(n6545), .B(n6544), .ZN(n6546)
         );
  AOI22_X1 U4833 ( .A1(n6588), .A2(mem_i_pc_o[8]), .B1(n6554), .B2(
        reset_vector_i[8]), .ZN(n6544) );
  NAND2_X1 U4834 ( .A1(n3319), .A2(csr_mepc_w[8]), .ZN(n6545) );
  AOI22_X1 U4835 ( .A1(mem_addr_w[29]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[29]), .ZN(n1459) );
  AOI22_X1 U4836 ( .A1(mem_addr_w[30]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[30]), .ZN(n1460) );
  AOI22_X1 U4837 ( .A1(mem_addr_w[31]), .A2(n4821), .B1(n4822), .B2(
        mem_d_addr_o[31]), .ZN(n1461) );
  AOI22_X1 U4838 ( .A1(n7990), .A2(n6410), .B1(n7987), .B2(n7992), .ZN(
        u_lsu_N16) );
  AOI22_X1 U4839 ( .A1(n7990), .A2(n6576), .B1(n7989), .B2(n7992), .ZN(
        add_x_67_B_3_) );
  AOI22_X1 U4840 ( .A1(n7990), .A2(n6573), .B1(n7991), .B2(n7992), .ZN(
        add_x_67_B_4_) );
  INV_X1 U4841 ( .A(n6543), .ZN(n2904) );
  AOI21_X1 U4842 ( .B1(U4_RSOP_173_C3_DATA1_12), .B2(n3363), .A(n6542), .ZN(
        n6543) );
  OAI211_X1 U4843 ( .C1(n6762), .C2(n6551), .A(n6541), .B(n6540), .ZN(n6542)
         );
  AOI22_X1 U4844 ( .A1(n6588), .A2(mem_i_pc_o[12]), .B1(n6554), .B2(
        reset_vector_i[12]), .ZN(n6540) );
  NAND2_X1 U4845 ( .A1(n3319), .A2(csr_mepc_w[12]), .ZN(n6541) );
  NAND4_X1 U4846 ( .A1(n6539), .A2(n6538), .A3(n6537), .A4(n6536), .ZN(n2903)
         );
  NAND2_X1 U4847 ( .A1(n6555), .A2(n_0_net__13_), .ZN(n6536) );
  NAND2_X1 U4848 ( .A1(n6589), .A2(csr_mepc_w[13]), .ZN(n6537) );
  AOI22_X1 U4849 ( .A1(n6588), .A2(mem_i_pc_o[13]), .B1(n6554), .B2(
        reset_vector_i[13]), .ZN(n6538) );
  NAND2_X1 U4850 ( .A1(U4_RSOP_173_C3_DATA1_13), .A2(n3363), .ZN(n6539) );
  INV_X1 U4851 ( .A(n6535), .ZN(n2900) );
  AOI21_X1 U4852 ( .B1(U4_RSOP_173_C3_DATA1_16), .B2(n3363), .A(n6534), .ZN(
        n6535) );
  OAI211_X1 U4853 ( .C1(n6763), .C2(n6551), .A(n6533), .B(n6532), .ZN(n6534)
         );
  AOI22_X1 U4854 ( .A1(n6588), .A2(mem_i_pc_o[16]), .B1(n6554), .B2(
        reset_vector_i[16]), .ZN(n6532) );
  NAND2_X1 U4855 ( .A1(n3319), .A2(csr_mepc_w[16]), .ZN(n6533) );
  NAND4_X1 U4856 ( .A1(n6531), .A2(n6530), .A3(n6529), .A4(n6528), .ZN(n2899)
         );
  NAND2_X1 U4857 ( .A1(n6555), .A2(n_0_net__17_), .ZN(n6528) );
  NAND2_X1 U4858 ( .A1(n3319), .A2(csr_mepc_w[17]), .ZN(n6529) );
  AOI22_X1 U4859 ( .A1(n6588), .A2(mem_i_pc_o[17]), .B1(n6554), .B2(
        reset_vector_i[17]), .ZN(n6530) );
  NAND2_X1 U4860 ( .A1(U4_RSOP_173_C3_DATA1_17), .A2(n3363), .ZN(n6531) );
  INV_X1 U4861 ( .A(exception_w), .ZN(n6683) );
  INV_X1 U4862 ( .A(n6527), .ZN(n2896) );
  AOI21_X1 U4863 ( .B1(U4_RSOP_173_C3_DATA1_20), .B2(n3363), .A(n6526), .ZN(
        n6527) );
  OAI211_X1 U4864 ( .C1(n6764), .C2(n6551), .A(n6525), .B(n6524), .ZN(n6526)
         );
  AOI22_X1 U4865 ( .A1(n6588), .A2(mem_i_pc_o[20]), .B1(n6554), .B2(
        reset_vector_i[20]), .ZN(n6524) );
  NAND2_X1 U4866 ( .A1(n3319), .A2(csr_mepc_w[20]), .ZN(n6525) );
  INV_X1 U4867 ( .A(n6523), .ZN(n2894) );
  AOI21_X1 U4868 ( .B1(U4_RSOP_173_C3_DATA1_22), .B2(n3363), .A(n6522), .ZN(
        n6523) );
  OAI211_X1 U4869 ( .C1(n6765), .C2(n6551), .A(n6521), .B(n6520), .ZN(n6522)
         );
  AOI22_X1 U4870 ( .A1(n6588), .A2(mem_i_pc_o[22]), .B1(n6554), .B2(
        reset_vector_i[22]), .ZN(n6520) );
  NAND2_X1 U4871 ( .A1(n3319), .A2(csr_mepc_w[22]), .ZN(n6521) );
  NAND4_X1 U4872 ( .A1(n6519), .A2(n6518), .A3(n6517), .A4(n6516), .ZN(n2893)
         );
  NAND2_X1 U4873 ( .A1(n6555), .A2(n_0_net__23_), .ZN(n6516) );
  NAND2_X1 U4874 ( .A1(n3319), .A2(csr_mepc_w[23]), .ZN(n6517) );
  AOI22_X1 U4875 ( .A1(n6588), .A2(mem_i_pc_o[23]), .B1(n6554), .B2(
        reset_vector_i[23]), .ZN(n6518) );
  NAND2_X1 U4876 ( .A1(U4_RSOP_173_C3_DATA1_23), .A2(n3363), .ZN(n6519) );
  INV_X1 U4877 ( .A(n6515), .ZN(n2892) );
  AOI21_X1 U4878 ( .B1(U4_RSOP_173_C3_DATA1_24), .B2(n3363), .A(n6514), .ZN(
        n6515) );
  OAI211_X1 U4879 ( .C1(n6766), .C2(n6551), .A(n6513), .B(n6512), .ZN(n6514)
         );
  AOI22_X1 U4880 ( .A1(n6588), .A2(mem_i_pc_o[24]), .B1(n6554), .B2(
        reset_vector_i[24]), .ZN(n6512) );
  NAND2_X1 U4881 ( .A1(n3319), .A2(csr_mepc_w[24]), .ZN(n6513) );
  NAND4_X1 U4882 ( .A1(n6511), .A2(n6510), .A3(n6509), .A4(n6508), .ZN(n2891)
         );
  NAND2_X1 U4883 ( .A1(n6555), .A2(n_0_net__25_), .ZN(n6508) );
  NOR2_X1 U4884 ( .A1(n6507), .A2(n6506), .ZN(n_0_net__25_) );
  AND2_X1 U4885 ( .A1(n6687), .A2(n6505), .ZN(n6506) );
  NAND2_X1 U4886 ( .A1(n3319), .A2(csr_mepc_w[25]), .ZN(n6509) );
  AOI22_X1 U4887 ( .A1(n6588), .A2(mem_i_pc_o[25]), .B1(n6554), .B2(
        reset_vector_i[25]), .ZN(n6510) );
  NAND2_X1 U4888 ( .A1(U4_RSOP_173_C3_DATA1_25), .A2(n3363), .ZN(n6511) );
  INV_X1 U4889 ( .A(n6504), .ZN(n2890) );
  AOI21_X1 U4890 ( .B1(U4_RSOP_173_C3_DATA1_26), .B2(n6559), .A(n6503), .ZN(
        n6504) );
  OAI211_X1 U4891 ( .C1(n6551), .C2(n6767), .A(n6502), .B(n6501), .ZN(n6503)
         );
  AOI22_X1 U4892 ( .A1(n6588), .A2(mem_i_pc_o[26]), .B1(n6554), .B2(
        reset_vector_i[26]), .ZN(n6501) );
  NAND2_X1 U4893 ( .A1(n3319), .A2(csr_mepc_w[26]), .ZN(n6502) );
  OAI21_X1 U4894 ( .B1(n6507), .B2(reset_vector_i[26]), .A(n6496), .ZN(n6767)
         );
  NAND4_X1 U4895 ( .A1(n6500), .A2(n6499), .A3(n6498), .A4(n6497), .ZN(n2889)
         );
  NAND2_X1 U4896 ( .A1(n_0_net__27_), .A2(n6555), .ZN(n6497) );
  AOI21_X1 U4897 ( .B1(n6496), .B2(n6495), .A(n6494), .ZN(n_0_net__27_) );
  NAND2_X1 U4898 ( .A1(n3319), .A2(csr_mepc_w[27]), .ZN(n6498) );
  AOI22_X1 U4899 ( .A1(n6588), .A2(mem_i_pc_o[27]), .B1(n6554), .B2(
        reset_vector_i[27]), .ZN(n6499) );
  NAND2_X1 U4900 ( .A1(U4_RSOP_173_C3_DATA1_27), .A2(n3363), .ZN(n6500) );
  OAI211_X1 U4901 ( .C1(n6551), .C2(n6768), .A(n6491), .B(n6490), .ZN(n2888)
         );
  AOI21_X1 U4902 ( .B1(n3319), .B2(csr_mepc_w[28]), .A(n6489), .ZN(n6490) );
  OAI22_X1 U4903 ( .A1(n6492), .A2(n3872), .B1(n6493), .B2(n6488), .ZN(n6489)
         );
  INV_X1 U4904 ( .A(reset_vector_i[28]), .ZN(n6488) );
  NAND2_X1 U4905 ( .A1(U4_RSOP_173_C3_DATA1_28), .A2(n3363), .ZN(n6491) );
  OAI21_X1 U4906 ( .B1(n6494), .B2(reset_vector_i[28]), .A(n6482), .ZN(n6768)
         );
  OAI211_X1 U4907 ( .C1(n6551), .C2(n6487), .A(n6486), .B(n6485), .ZN(n2887)
         );
  AOI21_X1 U4908 ( .B1(n3319), .B2(csr_mepc_w[29]), .A(n6484), .ZN(n6485) );
  OAI22_X1 U4909 ( .A1(n6492), .A2(n3871), .B1(n6493), .B2(n6483), .ZN(n6484)
         );
  NAND2_X1 U4910 ( .A1(U4_RSOP_173_C3_DATA1_29), .A2(n3363), .ZN(n6486) );
  INV_X1 U4911 ( .A(n_0_net__29_), .ZN(n6487) );
  AOI21_X1 U4912 ( .B1(n6482), .B2(n6483), .A(n6481), .ZN(n_0_net__29_) );
  OAI211_X1 U4913 ( .C1(n6551), .C2(n6769), .A(n6480), .B(n6479), .ZN(n2886)
         );
  AOI21_X1 U4914 ( .B1(n3319), .B2(csr_mepc_w[30]), .A(n6478), .ZN(n6479) );
  OAI22_X1 U4915 ( .A1(n6492), .A2(n3870), .B1(n6493), .B2(n6477), .ZN(n6478)
         );
  INV_X1 U4916 ( .A(reset_vector_i[30]), .ZN(n6477) );
  NAND2_X1 U4917 ( .A1(U4_RSOP_173_C3_DATA1_30), .A2(n3363), .ZN(n6480) );
  XNOR2_X1 U4918 ( .A(n6481), .B(reset_vector_i[30]), .ZN(n6769) );
  AOI21_X1 U4919 ( .B1(n3319), .B2(csr_mepc_w[31]), .A(n6475), .ZN(n6476) );
  OAI22_X1 U4920 ( .A1(n6492), .A2(n3869), .B1(n6493), .B2(n6474), .ZN(n6475)
         );
  NOR2_X1 U4921 ( .A1(n6760), .A2(rst_i), .ZN(n6493) );
  NAND2_X1 U4922 ( .A1(n6473), .A2(n6773), .ZN(n6492) );
  NAND2_X1 U4923 ( .A1(n6470), .A2(n6587), .ZN(n6471) );
  INV_X1 U4924 ( .A(n6469), .ZN(n6470) );
  OAI22_X1 U4925 ( .A1(n4819), .A2(n3869), .B1(n3345), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n121) );
  OAI21_X1 U4926 ( .B1(n6585), .B2(n7988), .A(n6584), .ZN(
        DP_OP_181_135_5161_n70) );
  OAI21_X1 U4927 ( .B1(n6586), .B2(n6583), .A(mem_i_inst_i[21]), .ZN(n6584) );
  OAI211_X1 U4928 ( .C1(n6585), .C2(n7987), .A(n6582), .B(n6581), .ZN(C1_Z_2)
         );
  OAI21_X1 U4929 ( .B1(n6586), .B2(n6583), .A(mem_i_inst_i[22]), .ZN(n6582) );
  INV_X1 U4930 ( .A(n6580), .ZN(DP_OP_181_135_5161_n72) );
  AOI21_X1 U4931 ( .B1(n3297), .B2(n6577), .A(n6576), .ZN(n6578) );
  INV_X1 U4932 ( .A(n6575), .ZN(DP_OP_181_135_5161_n73) );
  AOI21_X1 U4933 ( .B1(n3297), .B2(n6577), .A(n6573), .ZN(n6574) );
  OAI21_X1 U4934 ( .B1(n6585), .B2(n6824), .A(n6572), .ZN(
        DP_OP_181_135_5161_n74) );
  OAI21_X1 U4935 ( .B1(n6586), .B2(n6583), .A(mem_i_inst_i[25]), .ZN(n6572) );
  OAI21_X1 U4936 ( .B1(n6585), .B2(n6827), .A(n6571), .ZN(
        DP_OP_181_135_5161_n75) );
  OAI21_X1 U4937 ( .B1(n6586), .B2(n6583), .A(mem_i_inst_i[26]), .ZN(n6571) );
  OAI21_X1 U4938 ( .B1(n6585), .B2(n6830), .A(n6570), .ZN(
        DP_OP_181_135_5161_n76) );
  OAI21_X1 U4939 ( .B1(n6586), .B2(n6583), .A(mem_i_inst_i[27]), .ZN(n6570) );
  INV_X1 U4940 ( .A(n3523), .ZN(n6548) );
  INV_X1 U4941 ( .A(n6569), .ZN(DP_OP_181_135_5161_n77) );
  AOI21_X1 U4942 ( .B1(n3297), .B2(n6577), .A(n6567), .ZN(n6568) );
  OAI21_X1 U4943 ( .B1(n6585), .B2(n6566), .A(n6565), .ZN(
        DP_OP_181_135_5161_n78) );
  OAI21_X1 U4944 ( .B1(n6586), .B2(n6583), .A(mem_i_inst_i[29]), .ZN(n6565) );
  INV_X1 U4945 ( .A(mem_i_inst_i[29]), .ZN(n6566) );
  OAI22_X1 U4946 ( .A1(n4819), .A2(n3822), .B1(n3308), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n99) );
  OAI21_X1 U4947 ( .B1(n6585), .B2(n6564), .A(n6563), .ZN(
        DP_OP_181_135_5161_n79) );
  OAI21_X1 U4948 ( .B1(n6586), .B2(n6583), .A(mem_i_inst_i[30]), .ZN(n6563) );
  OAI22_X1 U4949 ( .A1(n4819), .A2(n3821), .B1(n3525), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n100) );
  AOI21_X1 U4950 ( .B1(n6583), .B2(mem_i_inst_i[20]), .A(n6561), .ZN(n6562) );
  OAI21_X1 U4951 ( .B1(n6685), .B2(n6577), .A(n6560), .ZN(
        DP_OP_181_135_5161_n81) );
  OAI22_X1 U4952 ( .A1(n4819), .A2(n3819), .B1(n3351), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n102) );
  OAI21_X1 U4953 ( .B1(n6684), .B2(n6577), .A(n6560), .ZN(
        DP_OP_181_135_5161_n82) );
  OAI22_X1 U4954 ( .A1(n3287), .A2(n3818), .B1(n3290), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n103) );
  OAI21_X1 U4955 ( .B1(n6821), .B2(n6577), .A(n6560), .ZN(
        DP_OP_181_135_5161_n83) );
  OAI22_X1 U4956 ( .A1(n4819), .A2(n3817), .B1(n3323), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n104) );
  OAI21_X1 U4957 ( .B1(n6604), .B2(n6577), .A(n6560), .ZN(
        DP_OP_181_135_5161_n84) );
  OAI22_X1 U4958 ( .A1(n3287), .A2(n3816), .B1(n3304), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n105) );
  OAI21_X1 U4959 ( .B1(n6608), .B2(n6577), .A(n6560), .ZN(
        DP_OP_181_135_5161_n85) );
  OAI22_X1 U4960 ( .A1(n4819), .A2(n3863), .B1(n3339), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n106) );
  OAI21_X1 U4961 ( .B1(n3520), .B2(n6577), .A(n6560), .ZN(
        DP_OP_181_135_5161_n86) );
  OAI22_X1 U4962 ( .A1(n3287), .A2(n3862), .B1(n3300), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n107) );
  OAI21_X1 U4963 ( .B1(n6615), .B2(n6577), .A(n6560), .ZN(
        DP_OP_181_135_5161_n87) );
  OAI22_X1 U4964 ( .A1(n4819), .A2(n3861), .B1(n3334), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n108) );
  OAI21_X1 U4965 ( .B1(n6619), .B2(n6577), .A(n6560), .ZN(
        DP_OP_181_135_5161_n88) );
  OAI22_X1 U4966 ( .A1(n3287), .A2(n3860), .B1(n3349), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n109) );
  OAI22_X1 U4967 ( .A1(n4819), .A2(n3859), .B1(n3341), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n110) );
  OAI22_X1 U4968 ( .A1(n3287), .A2(n3858), .B1(n3301), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n111) );
  OAI22_X1 U4969 ( .A1(n4819), .A2(n3857), .B1(n3344), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n112) );
  OAI22_X1 U4970 ( .A1(n3287), .A2(n3856), .B1(n3307), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n113) );
  OAI22_X1 U4971 ( .A1(n4819), .A2(n3855), .B1(n3335), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n114) );
  OAI22_X1 U4972 ( .A1(n3287), .A2(n3854), .B1(n3330), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n115) );
  OAI22_X1 U4973 ( .A1(n4819), .A2(n3853), .B1(n3333), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n116) );
  OAI22_X1 U4974 ( .A1(n3287), .A2(n3852), .B1(n3331), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n117) );
  OAI22_X1 U4975 ( .A1(n4819), .A2(n3872), .B1(n3320), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n118) );
  OAI22_X1 U4976 ( .A1(n4819), .A2(n3871), .B1(n3305), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n119) );
  NOR2_X1 U4977 ( .A1(n3297), .A2(n4910), .ZN(n6561) );
  OAI22_X1 U4978 ( .A1(n4819), .A2(n3870), .B1(n3347), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n120) );
  NAND2_X1 U4979 ( .A1(n4716), .A2(n4714), .ZN(n4713) );
  INV_X1 U4980 ( .A(n6742), .ZN(n4714) );
  INV_X1 U4981 ( .A(n4716), .ZN(n4715) );
  NOR2_X1 U4982 ( .A1(n6464), .A2(n4717), .ZN(n4716) );
  INV_X1 U4983 ( .A(n6458), .ZN(n4717) );
  AND2_X1 U4984 ( .A1(n6679), .A2(mem_i_inst_i[3]), .ZN(n6462) );
  NOR2_X1 U4985 ( .A1(n6461), .A2(n6679), .ZN(n6463) );
  NAND2_X1 U4986 ( .A1(n6460), .A2(n6469), .ZN(n6461) );
  NOR2_X1 U4987 ( .A1(n6457), .A2(mem_i_inst_i[3]), .ZN(n6458) );
  NAND2_X1 U4988 ( .A1(n6394), .A2(mem_i_inst_i[12]), .ZN(n6742) );
  INV_X1 U4989 ( .A(n6774), .ZN(n6394) );
  NAND2_X1 U4990 ( .A1(n6449), .A2(n6740), .ZN(n6448) );
  OAI211_X1 U4991 ( .C1(mem_i_inst_i[12]), .C2(u_branch_N125), .A(n6451), .B(
        n6680), .ZN(n6452) );
  OR2_X1 U4992 ( .A1(u_branch_N127), .A2(n6685), .ZN(n6451) );
  NAND4_X1 U4993 ( .A1(n6447), .A2(n3802), .A3(n3770), .A4(n6446), .ZN(n6449)
         );
  NOR2_X1 U4994 ( .A1(n6445), .A2(n6444), .ZN(n6446) );
  NAND3_X1 U4995 ( .A1(n6443), .A2(n6442), .A3(n6441), .ZN(n6444) );
  XNOR2_X1 U4996 ( .A(rs2_val_gpr_w[12]), .B(rs1_val_gpr_w[12]), .ZN(n6441) );
  AOI22_X1 U4997 ( .A1(n3346), .A2(rs1_val_gpr_w[30]), .B1(n3348), .B2(
        rs1_val_gpr_w[28]), .ZN(n6442) );
  AOI22_X1 U4998 ( .A1(n3339), .A2(rs2_val_gpr_w[16]), .B1(n3331), .B2(
        rs2_val_gpr_w[27]), .ZN(n6443) );
  NAND4_X1 U4999 ( .A1(n6440), .A2(n6439), .A3(n6438), .A4(n6437), .ZN(n6445)
         );
  AOI22_X1 U5000 ( .A1(n3304), .A2(rs2_val_gpr_w[15]), .B1(n3343), .B2(
        rs1_val_gpr_w[22]), .ZN(n6437) );
  AOI22_X1 U5001 ( .A1(n3330), .A2(rs2_val_gpr_w[25]), .B1(n3312), .B2(
        rs1_val_gpr_w[21]), .ZN(n6438) );
  AOI22_X1 U5002 ( .A1(n3289), .A2(rs2_val_gpr_w[11]), .B1(n3292), .B2(n3523), 
        .ZN(n6439) );
  AOI22_X1 U5003 ( .A1(n3321), .A2(rs2_val_gpr_w[8]), .B1(n3332), .B2(
        rs1_val_gpr_w[19]), .ZN(n6440) );
  AND4_X1 U5004 ( .A1(n6436), .A2(n6435), .A3(n6434), .A4(n6433), .ZN(n3770)
         );
  XNOR2_X1 U5005 ( .A(rs2_val_gpr_w[20]), .B(rs1_val_gpr_w[20]), .ZN(n6434) );
  XNOR2_X1 U5006 ( .A(rs2_val_gpr_w[3]), .B(rs1_val_gpr_w[3]), .ZN(n6435) );
  XNOR2_X1 U5007 ( .A(rs2_val_gpr_w[17]), .B(rs1_val_gpr_w[17]), .ZN(n6436) );
  AND4_X1 U5008 ( .A1(n6432), .A2(n6431), .A3(n6430), .A4(n6429), .ZN(n3802)
         );
  XNOR2_X1 U5009 ( .A(rs2_val_gpr_w[24]), .B(rs1_val_gpr_w[24]), .ZN(n6429) );
  XNOR2_X1 U5010 ( .A(rs2_val_gpr_w[5]), .B(rs1_val_gpr_w[5]), .ZN(n6431) );
  XNOR2_X1 U5011 ( .A(rs2_val_gpr_w[4]), .B(rs1_val_gpr_w[4]), .ZN(n6432) );
  NOR3_X1 U5012 ( .A1(n6428), .A2(n6427), .A3(n6426), .ZN(n6447) );
  NAND2_X1 U5013 ( .A1(n6425), .A2(n6424), .ZN(n6426) );
  XNOR2_X1 U5014 ( .A(rs2_val_gpr_w[29]), .B(rs1_val_gpr_w[29]), .ZN(n6424) );
  NAND4_X1 U5015 ( .A1(n6423), .A2(n6422), .A3(n6421), .A4(n6420), .ZN(n6428)
         );
  AOI21_X1 U5016 ( .B1(n3337), .B2(rs1_val_gpr_w[18]), .A(n6419), .ZN(n6420)
         );
  NAND3_X1 U5017 ( .A1(n6418), .A2(n6417), .A3(n6416), .ZN(n6419) );
  NOR2_X1 U5018 ( .A1(n6731), .A2(n6730), .ZN(n6416) );
  NOR4_X1 U5019 ( .A1(n6739), .A2(n6738), .A3(n6737), .A4(n6736), .ZN(n6417)
         );
  NOR4_X1 U5020 ( .A1(n6735), .A2(n6734), .A3(n6733), .A4(n6732), .ZN(n6418)
         );
  AOI22_X1 U5021 ( .A1(n3323), .A2(rs2_val_gpr_w[14]), .B1(n3313), .B2(
        rs1_val_gpr_w[6]), .ZN(n6421) );
  AOI22_X1 U5022 ( .A1(n3308), .A2(rs2_val_gpr_w[9]), .B1(n3291), .B2(
        rs1_val_gpr_w[13]), .ZN(n6422) );
  AOI22_X1 U5023 ( .A1(n3333), .A2(rs2_val_gpr_w[26]), .B1(n3307), .B2(
        rs2_val_gpr_w[23]), .ZN(n6423) );
  INV_X1 U5024 ( .A(n6681), .ZN(n6450) );
  INV_X1 U5025 ( .A(n6682), .ZN(n6455) );
  NOR2_X1 U5026 ( .A1(n6774), .A2(mem_i_inst_i[12]), .ZN(n6682) );
  NAND2_X1 U5027 ( .A1(n6684), .A2(mem_i_inst_i[14]), .ZN(n6774) );
  NAND2_X1 U5028 ( .A1(n3298), .A2(rs1_val_gpr_w[31]), .ZN(n6741) );
  NAND2_X1 U5029 ( .A1(n3345), .A2(rs2_val_gpr_w[31]), .ZN(n6740) );
  AOI22_X1 U5030 ( .A1(reg_file[799]), .A2(n4788), .B1(n4787), .B2(
        reg_file[831]), .ZN(n5814) );
  AOI22_X1 U5031 ( .A1(reg_file[895]), .A2(n4778), .B1(n3799), .B2(
        reg_file[863]), .ZN(n5815) );
  AOI22_X1 U5032 ( .A1(n4818), .A2(reg_file[959]), .B1(n3769), .B2(
        reg_file[927]), .ZN(n5816) );
  AOI22_X1 U5033 ( .A1(reg_file[1023]), .A2(n4758), .B1(n4757), .B2(
        reg_file[991]), .ZN(n5817) );
  AOI22_X1 U5034 ( .A1(reg_file[639]), .A2(n4778), .B1(n3799), .B2(
        reg_file[607]), .ZN(n5806) );
  AOI22_X1 U5035 ( .A1(n4818), .A2(reg_file[703]), .B1(n3769), .B2(
        reg_file[671]), .ZN(n5807) );
  AOI22_X1 U5036 ( .A1(n4812), .A2(reg_file[543]), .B1(n4809), .B2(
        reg_file[575]), .ZN(n6388) );
  AOI22_X1 U5037 ( .A1(n3285), .A2(reg_file[639]), .B1(n4806), .B2(
        reg_file[607]), .ZN(n6389) );
  AOI22_X1 U5038 ( .A1(n4801), .A2(reg_file[735]), .B1(n4797), .B2(
        reg_file[703]), .ZN(n6390) );
  AOI22_X1 U5039 ( .A1(n3355), .A2(reg_file[671]), .B1(n4813), .B2(
        reg_file[767]), .ZN(n6391) );
  AOI22_X1 U5040 ( .A1(n3286), .A2(reg_file[383]), .B1(n4806), .B2(
        reg_file[351]), .ZN(n6378) );
  AOI22_X1 U5041 ( .A1(n4801), .A2(reg_file[479]), .B1(n4797), .B2(
        reg_file[447]), .ZN(n6379) );
  AOI22_X1 U5042 ( .A1(n3386), .A2(reg_file[415]), .B1(n3293), .B2(
        reg_file[511]), .ZN(n6380) );
  AOI22_X1 U5043 ( .A1(n4812), .A2(reg_file[799]), .B1(n4809), .B2(
        reg_file[831]), .ZN(n6374) );
  AOI22_X1 U5044 ( .A1(n3285), .A2(reg_file[895]), .B1(n4806), .B2(
        reg_file[863]), .ZN(n6375) );
  AOI22_X1 U5045 ( .A1(n4801), .A2(reg_file[991]), .B1(n4797), .B2(
        reg_file[959]), .ZN(n6376) );
  AOI22_X1 U5046 ( .A1(n3355), .A2(reg_file[927]), .B1(n4814), .B2(
        reg_file[1023]), .ZN(n6377) );
  AOI22_X1 U5047 ( .A1(n4811), .A2(reg_file[31]), .B1(n4809), .B2(reg_file[63]), .ZN(n6369) );
  AOI22_X1 U5048 ( .A1(n3286), .A2(reg_file[127]), .B1(n4806), .B2(
        reg_file[95]), .ZN(n6370) );
  AOI22_X1 U5049 ( .A1(n4801), .A2(reg_file[223]), .B1(n4797), .B2(
        reg_file[191]), .ZN(n6371) );
  AOI22_X1 U5050 ( .A1(n3355), .A2(reg_file[159]), .B1(n4813), .B2(
        reg_file[255]), .ZN(n6372) );
  NAND2_X1 U5051 ( .A1(n6224), .A2(n3362), .ZN(n6225) );
  NAND4_X1 U5052 ( .A1(n6223), .A2(n6222), .A3(n6221), .A4(n6220), .ZN(n6224)
         );
  AOI22_X1 U5053 ( .A1(n3358), .A2(reg_file[786]), .B1(n4809), .B2(
        reg_file[818]), .ZN(n6220) );
  AOI22_X1 U5054 ( .A1(n3285), .A2(reg_file[882]), .B1(n3359), .B2(
        reg_file[850]), .ZN(n6221) );
  AOI22_X1 U5055 ( .A1(n3356), .A2(reg_file[978]), .B1(n3360), .B2(
        reg_file[946]), .ZN(n6222) );
  AOI22_X1 U5056 ( .A1(n3355), .A2(reg_file[914]), .B1(n4813), .B2(
        reg_file[1010]), .ZN(n6223) );
  NAND2_X1 U5057 ( .A1(n6219), .A2(n3387), .ZN(n6226) );
  NAND4_X1 U5058 ( .A1(n6218), .A2(n6217), .A3(n6216), .A4(n6215), .ZN(n6219)
         );
  AOI22_X1 U5059 ( .A1(n3358), .A2(reg_file[274]), .B1(n4809), .B2(
        reg_file[306]), .ZN(n6215) );
  AOI22_X1 U5060 ( .A1(n3286), .A2(reg_file[370]), .B1(n3359), .B2(
        reg_file[338]), .ZN(n6216) );
  AOI22_X1 U5061 ( .A1(n3356), .A2(reg_file[466]), .B1(n3360), .B2(
        reg_file[434]), .ZN(n6217) );
  AOI22_X1 U5062 ( .A1(n3355), .A2(reg_file[402]), .B1(n4813), .B2(
        reg_file[498]), .ZN(n6218) );
  NAND2_X1 U5063 ( .A1(n6214), .A2(n3388), .ZN(n6227) );
  NAND4_X1 U5064 ( .A1(n6213), .A2(n6212), .A3(n6211), .A4(n6210), .ZN(n6214)
         );
  AOI22_X1 U5065 ( .A1(n3358), .A2(reg_file[530]), .B1(n4809), .B2(
        reg_file[562]), .ZN(n6210) );
  AOI22_X1 U5066 ( .A1(n3285), .A2(reg_file[626]), .B1(n3359), .B2(
        reg_file[594]), .ZN(n6211) );
  AOI22_X1 U5067 ( .A1(n3356), .A2(reg_file[722]), .B1(n3360), .B2(
        reg_file[690]), .ZN(n6212) );
  AOI22_X1 U5068 ( .A1(n3355), .A2(reg_file[658]), .B1(n4813), .B2(
        reg_file[754]), .ZN(n6213) );
  NAND2_X1 U5069 ( .A1(n6209), .A2(n6373), .ZN(n6228) );
  NAND4_X1 U5070 ( .A1(n6208), .A2(n6207), .A3(n6206), .A4(n6205), .ZN(n6209)
         );
  AOI22_X1 U5071 ( .A1(n3358), .A2(reg_file[18]), .B1(n4809), .B2(reg_file[50]), .ZN(n6205) );
  AOI22_X1 U5072 ( .A1(n3286), .A2(reg_file[114]), .B1(n3359), .B2(
        reg_file[82]), .ZN(n6206) );
  AOI22_X1 U5073 ( .A1(n3356), .A2(reg_file[210]), .B1(n3360), .B2(
        reg_file[178]), .ZN(n6207) );
  AOI22_X1 U5074 ( .A1(n3386), .A2(reg_file[146]), .B1(n4813), .B2(
        reg_file[242]), .ZN(n6208) );
  NAND4_X1 U5075 ( .A1(n5539), .A2(n5538), .A3(n5537), .A4(n5536), .ZN(
        rs2_val_gpr_w[18]) );
  NAND2_X1 U5076 ( .A1(n5535), .A2(n3390), .ZN(n5536) );
  NAND4_X1 U5077 ( .A1(n5534), .A2(n5533), .A3(n5532), .A4(n5531), .ZN(n5535)
         );
  AOI22_X1 U5078 ( .A1(n4788), .A2(reg_file[530]), .B1(n4786), .B2(
        reg_file[562]), .ZN(n5531) );
  AOI22_X1 U5079 ( .A1(n4782), .A2(reg_file[626]), .B1(n4775), .B2(
        reg_file[594]), .ZN(n5532) );
  AOI22_X1 U5080 ( .A1(n3294), .A2(reg_file[690]), .B1(n4766), .B2(
        reg_file[658]), .ZN(n5533) );
  AOI22_X1 U5081 ( .A1(n4757), .A2(reg_file[722]), .B1(n4758), .B2(
        reg_file[754]), .ZN(n5534) );
  NAND2_X1 U5082 ( .A1(n5530), .A2(n3389), .ZN(n5537) );
  NAND4_X1 U5083 ( .A1(n5529), .A2(n5528), .A3(n5527), .A4(n5526), .ZN(n5530)
         );
  AOI22_X1 U5084 ( .A1(n4788), .A2(reg_file[274]), .B1(n4786), .B2(
        reg_file[306]), .ZN(n5526) );
  AOI22_X1 U5085 ( .A1(n4782), .A2(reg_file[370]), .B1(n4775), .B2(
        reg_file[338]), .ZN(n5527) );
  AOI22_X1 U5086 ( .A1(n3294), .A2(reg_file[434]), .B1(n4766), .B2(
        reg_file[402]), .ZN(n5528) );
  AOI22_X1 U5087 ( .A1(n4755), .A2(reg_file[466]), .B1(n4758), .B2(
        reg_file[498]), .ZN(n5529) );
  NAND2_X1 U5088 ( .A1(n5525), .A2(n3361), .ZN(n5538) );
  NAND4_X1 U5089 ( .A1(n5524), .A2(n5523), .A3(n5522), .A4(n5521), .ZN(n5525)
         );
  AOI22_X1 U5090 ( .A1(n4788), .A2(reg_file[786]), .B1(n4786), .B2(
        reg_file[818]), .ZN(n5521) );
  AOI22_X1 U5091 ( .A1(n4782), .A2(reg_file[882]), .B1(n4775), .B2(
        reg_file[850]), .ZN(n5522) );
  AOI22_X1 U5092 ( .A1(n3294), .A2(reg_file[946]), .B1(n4766), .B2(
        reg_file[914]), .ZN(n5523) );
  AOI22_X1 U5093 ( .A1(n5809), .A2(reg_file[978]), .B1(n4758), .B2(
        reg_file[1010]), .ZN(n5524) );
  NAND2_X1 U5094 ( .A1(n5520), .A2(n4754), .ZN(n5539) );
  NAND4_X1 U5095 ( .A1(n5519), .A2(n5518), .A3(n5517), .A4(n5516), .ZN(n5520)
         );
  AOI22_X1 U5096 ( .A1(n4788), .A2(reg_file[18]), .B1(n4786), .B2(reg_file[50]), .ZN(n5516) );
  AOI22_X1 U5097 ( .A1(n4782), .A2(reg_file[114]), .B1(n4775), .B2(
        reg_file[82]), .ZN(n5517) );
  AOI22_X1 U5098 ( .A1(n3294), .A2(reg_file[178]), .B1(n4766), .B2(
        reg_file[146]), .ZN(n5518) );
  AOI22_X1 U5099 ( .A1(n4757), .A2(reg_file[210]), .B1(n4758), .B2(
        reg_file[242]), .ZN(n5519) );
  NAND4_X1 U5100 ( .A1(n6245), .A2(n6244), .A3(n6243), .A4(n6242), .ZN(n6246)
         );
  AOI22_X1 U5101 ( .A1(n3358), .A2(reg_file[531]), .B1(n4809), .B2(
        reg_file[563]), .ZN(n6242) );
  AOI22_X1 U5102 ( .A1(n3285), .A2(reg_file[627]), .B1(n3359), .B2(
        reg_file[595]), .ZN(n6243) );
  AOI22_X1 U5103 ( .A1(n3356), .A2(reg_file[723]), .B1(n3360), .B2(
        reg_file[691]), .ZN(n6244) );
  AOI22_X1 U5104 ( .A1(n3355), .A2(reg_file[659]), .B1(n4815), .B2(
        reg_file[755]), .ZN(n6245) );
  NAND4_X1 U5105 ( .A1(n6240), .A2(n6239), .A3(n6238), .A4(n6237), .ZN(n6241)
         );
  AOI22_X1 U5106 ( .A1(n3358), .A2(reg_file[19]), .B1(n4809), .B2(reg_file[51]), .ZN(n6237) );
  AOI22_X1 U5107 ( .A1(n3285), .A2(reg_file[115]), .B1(n3359), .B2(
        reg_file[83]), .ZN(n6238) );
  AOI22_X1 U5108 ( .A1(n3356), .A2(reg_file[211]), .B1(n3360), .B2(
        reg_file[179]), .ZN(n6239) );
  AOI22_X1 U5109 ( .A1(n3386), .A2(reg_file[147]), .B1(n4813), .B2(
        reg_file[243]), .ZN(n6240) );
  AOI22_X1 U5110 ( .A1(n3358), .A2(reg_file[787]), .B1(n4809), .B2(
        reg_file[819]), .ZN(n6233) );
  AOI22_X1 U5111 ( .A1(n3286), .A2(reg_file[883]), .B1(n3359), .B2(
        reg_file[851]), .ZN(n6234) );
  AOI22_X1 U5112 ( .A1(n3356), .A2(reg_file[979]), .B1(n3360), .B2(
        reg_file[947]), .ZN(n6235) );
  AOI22_X1 U5113 ( .A1(n3355), .A2(reg_file[915]), .B1(n4815), .B2(
        reg_file[1011]), .ZN(n6236) );
  AOI22_X1 U5114 ( .A1(n3358), .A2(reg_file[275]), .B1(n4809), .B2(
        reg_file[307]), .ZN(n6229) );
  AOI22_X1 U5115 ( .A1(n3285), .A2(reg_file[371]), .B1(n3359), .B2(
        reg_file[339]), .ZN(n6230) );
  AOI22_X1 U5116 ( .A1(n3356), .A2(reg_file[467]), .B1(n3360), .B2(
        reg_file[435]), .ZN(n6231) );
  AOI22_X1 U5117 ( .A1(n3355), .A2(reg_file[403]), .B1(n4815), .B2(
        reg_file[499]), .ZN(n6232) );
  NAND4_X1 U5118 ( .A1(n5563), .A2(n5562), .A3(n5561), .A4(n5560), .ZN(
        rs2_val_gpr_w[19]) );
  NAND2_X1 U5119 ( .A1(n5559), .A2(n3361), .ZN(n5560) );
  NAND4_X1 U5120 ( .A1(n5558), .A2(n5557), .A3(n5556), .A4(n5555), .ZN(n5559)
         );
  AOI22_X1 U5121 ( .A1(n4788), .A2(reg_file[787]), .B1(n4786), .B2(
        reg_file[819]), .ZN(n5555) );
  AOI22_X1 U5122 ( .A1(n4781), .A2(reg_file[883]), .B1(n4775), .B2(
        reg_file[851]), .ZN(n5556) );
  AOI22_X1 U5123 ( .A1(n3294), .A2(reg_file[947]), .B1(n4766), .B2(
        reg_file[915]), .ZN(n5557) );
  AOI22_X1 U5124 ( .A1(n4757), .A2(reg_file[979]), .B1(n4758), .B2(
        reg_file[1011]), .ZN(n5558) );
  NAND2_X1 U5125 ( .A1(n5554), .A2(n3390), .ZN(n5561) );
  NAND4_X1 U5126 ( .A1(n5553), .A2(n5552), .A3(n5551), .A4(n5550), .ZN(n5554)
         );
  AOI22_X1 U5127 ( .A1(n4788), .A2(reg_file[531]), .B1(n4786), .B2(
        reg_file[563]), .ZN(n5550) );
  AOI22_X1 U5128 ( .A1(n4781), .A2(reg_file[627]), .B1(n4775), .B2(
        reg_file[595]), .ZN(n5551) );
  AOI22_X1 U5129 ( .A1(n3294), .A2(reg_file[691]), .B1(n4766), .B2(
        reg_file[659]), .ZN(n5552) );
  AOI22_X1 U5130 ( .A1(n3519), .A2(reg_file[723]), .B1(n4758), .B2(
        reg_file[755]), .ZN(n5553) );
  NAND2_X1 U5131 ( .A1(n5549), .A2(n4754), .ZN(n5562) );
  NAND4_X1 U5132 ( .A1(n5548), .A2(n5547), .A3(n5546), .A4(n5545), .ZN(n5549)
         );
  AOI22_X1 U5133 ( .A1(n4788), .A2(reg_file[19]), .B1(n4786), .B2(reg_file[51]), .ZN(n5545) );
  AOI22_X1 U5134 ( .A1(n4781), .A2(reg_file[115]), .B1(n4775), .B2(
        reg_file[83]), .ZN(n5546) );
  AOI22_X1 U5135 ( .A1(n3294), .A2(reg_file[179]), .B1(n4766), .B2(
        reg_file[147]), .ZN(n5547) );
  AOI22_X1 U5136 ( .A1(n4757), .A2(reg_file[211]), .B1(n4758), .B2(
        reg_file[243]), .ZN(n5548) );
  NAND2_X1 U5137 ( .A1(n5544), .A2(n3389), .ZN(n5563) );
  NAND4_X1 U5138 ( .A1(n5543), .A2(n5542), .A3(n5541), .A4(n5540), .ZN(n5544)
         );
  AOI22_X1 U5139 ( .A1(n4788), .A2(reg_file[275]), .B1(n4786), .B2(
        reg_file[307]), .ZN(n5540) );
  AOI22_X1 U5140 ( .A1(n4781), .A2(reg_file[371]), .B1(n4775), .B2(
        reg_file[339]), .ZN(n5541) );
  AOI22_X1 U5141 ( .A1(n3294), .A2(reg_file[435]), .B1(n4766), .B2(
        reg_file[403]), .ZN(n5542) );
  AOI22_X1 U5142 ( .A1(n4757), .A2(reg_file[467]), .B1(n4758), .B2(
        reg_file[499]), .ZN(n5543) );
  NAND4_X1 U5143 ( .A1(n6264), .A2(n6263), .A3(n6262), .A4(n6261), .ZN(n6265)
         );
  AOI22_X1 U5144 ( .A1(n3358), .A2(reg_file[788]), .B1(n4809), .B2(
        reg_file[820]), .ZN(n6261) );
  AOI22_X1 U5145 ( .A1(n3285), .A2(reg_file[884]), .B1(n3359), .B2(
        reg_file[852]), .ZN(n6262) );
  AOI22_X1 U5146 ( .A1(n3356), .A2(reg_file[980]), .B1(n3360), .B2(
        reg_file[948]), .ZN(n6263) );
  AOI22_X1 U5147 ( .A1(n3355), .A2(reg_file[916]), .B1(n4813), .B2(
        reg_file[1012]), .ZN(n6264) );
  NAND4_X1 U5148 ( .A1(n6259), .A2(n6258), .A3(n6257), .A4(n6256), .ZN(n6260)
         );
  AOI22_X1 U5149 ( .A1(n3358), .A2(reg_file[276]), .B1(n4809), .B2(
        reg_file[308]), .ZN(n6256) );
  AOI22_X1 U5150 ( .A1(n3286), .A2(reg_file[372]), .B1(n3359), .B2(
        reg_file[340]), .ZN(n6257) );
  AOI22_X1 U5151 ( .A1(n3356), .A2(reg_file[468]), .B1(n3360), .B2(
        reg_file[436]), .ZN(n6258) );
  AOI22_X1 U5152 ( .A1(n3355), .A2(reg_file[404]), .B1(n4813), .B2(
        reg_file[500]), .ZN(n6259) );
  NAND4_X1 U5153 ( .A1(n6254), .A2(n6253), .A3(n6252), .A4(n6251), .ZN(n6255)
         );
  AOI22_X1 U5154 ( .A1(n3358), .A2(reg_file[532]), .B1(n4809), .B2(
        reg_file[564]), .ZN(n6251) );
  AOI22_X1 U5155 ( .A1(n3285), .A2(reg_file[628]), .B1(n3359), .B2(
        reg_file[596]), .ZN(n6252) );
  AOI22_X1 U5156 ( .A1(n3356), .A2(reg_file[724]), .B1(n3360), .B2(
        reg_file[692]), .ZN(n6253) );
  AOI22_X1 U5157 ( .A1(n4790), .A2(reg_file[660]), .B1(n4813), .B2(
        reg_file[756]), .ZN(n6254) );
  AOI22_X1 U5158 ( .A1(n3358), .A2(reg_file[20]), .B1(n4809), .B2(reg_file[52]), .ZN(n6247) );
  AOI22_X1 U5159 ( .A1(n3286), .A2(reg_file[116]), .B1(n3359), .B2(
        reg_file[84]), .ZN(n6248) );
  AOI22_X1 U5160 ( .A1(n3356), .A2(reg_file[212]), .B1(n3360), .B2(
        reg_file[180]), .ZN(n6249) );
  AOI22_X1 U5161 ( .A1(n3355), .A2(reg_file[148]), .B1(n4813), .B2(
        reg_file[244]), .ZN(n6250) );
  NAND4_X1 U5162 ( .A1(n5587), .A2(n5586), .A3(n5585), .A4(n5584), .ZN(
        rs2_val_gpr_w[20]) );
  NAND2_X1 U5163 ( .A1(n5583), .A2(n3361), .ZN(n5584) );
  NAND4_X1 U5164 ( .A1(n5582), .A2(n5581), .A3(n5580), .A4(n5579), .ZN(n5583)
         );
  AOI22_X1 U5165 ( .A1(n4788), .A2(reg_file[788]), .B1(n4786), .B2(
        reg_file[820]), .ZN(n5579) );
  AOI22_X1 U5166 ( .A1(n4781), .A2(reg_file[884]), .B1(n4775), .B2(
        reg_file[852]), .ZN(n5580) );
  AOI22_X1 U5167 ( .A1(n3294), .A2(reg_file[948]), .B1(n4766), .B2(
        reg_file[916]), .ZN(n5581) );
  AOI22_X1 U5168 ( .A1(n4757), .A2(reg_file[980]), .B1(n4758), .B2(
        reg_file[1012]), .ZN(n5582) );
  NAND2_X1 U5169 ( .A1(n5578), .A2(n3389), .ZN(n5585) );
  NAND4_X1 U5170 ( .A1(n5577), .A2(n5576), .A3(n5575), .A4(n5574), .ZN(n5578)
         );
  AOI22_X1 U5171 ( .A1(n4788), .A2(reg_file[276]), .B1(n4786), .B2(
        reg_file[308]), .ZN(n5574) );
  AOI22_X1 U5172 ( .A1(n4781), .A2(reg_file[372]), .B1(n4775), .B2(
        reg_file[340]), .ZN(n5575) );
  AOI22_X1 U5173 ( .A1(n3294), .A2(reg_file[436]), .B1(n4766), .B2(
        reg_file[404]), .ZN(n5576) );
  AOI22_X1 U5174 ( .A1(n4757), .A2(reg_file[468]), .B1(n4758), .B2(
        reg_file[500]), .ZN(n5577) );
  NAND2_X1 U5175 ( .A1(n5573), .A2(n3390), .ZN(n5586) );
  NAND4_X1 U5176 ( .A1(n5572), .A2(n5571), .A3(n5570), .A4(n5569), .ZN(n5573)
         );
  AOI22_X1 U5177 ( .A1(n4788), .A2(reg_file[532]), .B1(n4786), .B2(
        reg_file[564]), .ZN(n5569) );
  AOI22_X1 U5178 ( .A1(n4781), .A2(reg_file[628]), .B1(n4775), .B2(
        reg_file[596]), .ZN(n5570) );
  AOI22_X1 U5179 ( .A1(n3294), .A2(reg_file[692]), .B1(n4766), .B2(
        reg_file[660]), .ZN(n5571) );
  AOI22_X1 U5180 ( .A1(n4757), .A2(reg_file[724]), .B1(n4758), .B2(
        reg_file[756]), .ZN(n5572) );
  NAND2_X1 U5181 ( .A1(n5568), .A2(n4754), .ZN(n5587) );
  NAND4_X1 U5182 ( .A1(n5567), .A2(n5566), .A3(n5565), .A4(n5564), .ZN(n5568)
         );
  AOI22_X1 U5183 ( .A1(n4788), .A2(reg_file[20]), .B1(n4786), .B2(reg_file[52]), .ZN(n5564) );
  AOI22_X1 U5184 ( .A1(n4781), .A2(reg_file[116]), .B1(n4775), .B2(
        reg_file[84]), .ZN(n5565) );
  BUF_X1 U5185 ( .A(n3799), .Z(n4775) );
  AOI22_X1 U5186 ( .A1(n3294), .A2(reg_file[180]), .B1(n4766), .B2(
        reg_file[148]), .ZN(n5566) );
  AOI22_X1 U5187 ( .A1(n4756), .A2(reg_file[212]), .B1(n4758), .B2(
        reg_file[244]), .ZN(n5567) );
  AOI22_X1 U5188 ( .A1(n3358), .A2(reg_file[789]), .B1(n4809), .B2(
        reg_file[821]), .ZN(n6270) );
  AOI22_X1 U5189 ( .A1(n3285), .A2(reg_file[885]), .B1(n3359), .B2(
        reg_file[853]), .ZN(n6271) );
  AOI22_X1 U5190 ( .A1(n3356), .A2(reg_file[981]), .B1(n4795), .B2(
        reg_file[949]), .ZN(n6272) );
  AOI22_X1 U5191 ( .A1(n3355), .A2(reg_file[917]), .B1(n3354), .B2(
        reg_file[1013]), .ZN(n6273) );
  AOI22_X1 U5192 ( .A1(n3358), .A2(reg_file[21]), .B1(n4808), .B2(reg_file[53]), .ZN(n6266) );
  AOI22_X1 U5193 ( .A1(n3286), .A2(reg_file[117]), .B1(n3359), .B2(
        reg_file[85]), .ZN(n6267) );
  AOI22_X1 U5194 ( .A1(n3356), .A2(reg_file[213]), .B1(n4795), .B2(
        reg_file[181]), .ZN(n6268) );
  AOI22_X1 U5195 ( .A1(n3355), .A2(reg_file[149]), .B1(n4815), .B2(
        reg_file[245]), .ZN(n6269) );
  NAND4_X1 U5196 ( .A1(n5611), .A2(n5610), .A3(n5609), .A4(n5608), .ZN(
        rs2_val_gpr_w[21]) );
  NAND2_X1 U5197 ( .A1(n5607), .A2(n3361), .ZN(n5608) );
  NAND4_X1 U5198 ( .A1(n5606), .A2(n5605), .A3(n5604), .A4(n5603), .ZN(n5607)
         );
  AOI22_X1 U5199 ( .A1(n4788), .A2(reg_file[789]), .B1(n4786), .B2(
        reg_file[821]), .ZN(n5603) );
  AOI22_X1 U5200 ( .A1(n4781), .A2(reg_file[885]), .B1(n4776), .B2(
        reg_file[853]), .ZN(n5604) );
  AOI22_X1 U5201 ( .A1(n3294), .A2(reg_file[949]), .B1(n3769), .B2(
        reg_file[917]), .ZN(n5605) );
  AOI22_X1 U5202 ( .A1(n4757), .A2(reg_file[981]), .B1(n4758), .B2(
        reg_file[1013]), .ZN(n5606) );
  NAND2_X1 U5203 ( .A1(n5602), .A2(n4754), .ZN(n5609) );
  NAND4_X1 U5204 ( .A1(n5601), .A2(n5600), .A3(n5599), .A4(n5598), .ZN(n5602)
         );
  AOI22_X1 U5205 ( .A1(n4788), .A2(reg_file[21]), .B1(n4787), .B2(reg_file[53]), .ZN(n5598) );
  AOI22_X1 U5206 ( .A1(n4781), .A2(reg_file[117]), .B1(n4776), .B2(
        reg_file[85]), .ZN(n5599) );
  AOI22_X1 U5207 ( .A1(n3294), .A2(reg_file[181]), .B1(n3769), .B2(
        reg_file[149]), .ZN(n5600) );
  AOI22_X1 U5208 ( .A1(n4757), .A2(reg_file[213]), .B1(n4758), .B2(
        reg_file[245]), .ZN(n5601) );
  NAND2_X1 U5209 ( .A1(n5597), .A2(n3390), .ZN(n5610) );
  NAND4_X1 U5210 ( .A1(n5596), .A2(n5595), .A3(n5594), .A4(n5593), .ZN(n5597)
         );
  AOI22_X1 U5211 ( .A1(n4788), .A2(reg_file[533]), .B1(n4787), .B2(
        reg_file[565]), .ZN(n5593) );
  AOI22_X1 U5212 ( .A1(n4781), .A2(reg_file[629]), .B1(n4776), .B2(
        reg_file[597]), .ZN(n5594) );
  AOI22_X1 U5213 ( .A1(n3294), .A2(reg_file[693]), .B1(n3769), .B2(
        reg_file[661]), .ZN(n5595) );
  AOI22_X1 U5214 ( .A1(n4755), .A2(reg_file[725]), .B1(n4758), .B2(
        reg_file[757]), .ZN(n5596) );
  NAND2_X1 U5215 ( .A1(n5592), .A2(n3389), .ZN(n5611) );
  NAND4_X1 U5216 ( .A1(n5591), .A2(n5590), .A3(n5589), .A4(n5588), .ZN(n5592)
         );
  AOI22_X1 U5217 ( .A1(n4788), .A2(reg_file[277]), .B1(n4786), .B2(
        reg_file[309]), .ZN(n5588) );
  AOI22_X1 U5218 ( .A1(n4781), .A2(reg_file[373]), .B1(n4776), .B2(
        reg_file[341]), .ZN(n5589) );
  AOI22_X1 U5219 ( .A1(n3294), .A2(reg_file[437]), .B1(n3769), .B2(
        reg_file[405]), .ZN(n5590) );
  AOI22_X1 U5220 ( .A1(n4756), .A2(reg_file[469]), .B1(n4758), .B2(
        reg_file[501]), .ZN(n5591) );
  NAND2_X1 U5221 ( .A1(n6200), .A2(n3362), .ZN(n6201) );
  NAND4_X1 U5222 ( .A1(n6199), .A2(n6198), .A3(n6197), .A4(n6196), .ZN(n6200)
         );
  AOI22_X1 U5223 ( .A1(n3316), .A2(reg_file[785]), .B1(n3315), .B2(
        reg_file[817]), .ZN(n6196) );
  AOI22_X1 U5224 ( .A1(n3314), .A2(reg_file[977]), .B1(n4794), .B2(
        reg_file[945]), .ZN(n6198) );
  AOI22_X1 U5225 ( .A1(n3386), .A2(reg_file[913]), .B1(n4813), .B2(
        reg_file[1009]), .ZN(n6199) );
  NAND2_X1 U5226 ( .A1(n6195), .A2(n3387), .ZN(n6202) );
  NAND4_X1 U5227 ( .A1(n6194), .A2(n6193), .A3(n6192), .A4(n6191), .ZN(n6195)
         );
  AOI22_X1 U5228 ( .A1(n3316), .A2(reg_file[273]), .B1(n3315), .B2(
        reg_file[305]), .ZN(n6191) );
  AOI22_X1 U5229 ( .A1(n3286), .A2(reg_file[369]), .B1(n4805), .B2(
        reg_file[337]), .ZN(n6192) );
  AOI22_X1 U5230 ( .A1(n3314), .A2(reg_file[465]), .B1(n4794), .B2(
        reg_file[433]), .ZN(n6193) );
  AOI22_X1 U5231 ( .A1(n3355), .A2(reg_file[401]), .B1(n4813), .B2(
        reg_file[497]), .ZN(n6194) );
  NAND2_X1 U5232 ( .A1(n6190), .A2(n3388), .ZN(n6203) );
  NAND4_X1 U5233 ( .A1(n6189), .A2(n6188), .A3(n6187), .A4(n6186), .ZN(n6190)
         );
  AOI22_X1 U5234 ( .A1(n3316), .A2(reg_file[529]), .B1(n3315), .B2(
        reg_file[561]), .ZN(n6186) );
  AOI22_X1 U5235 ( .A1(n3285), .A2(reg_file[625]), .B1(n4806), .B2(
        reg_file[593]), .ZN(n6187) );
  AOI22_X1 U5236 ( .A1(n3314), .A2(reg_file[721]), .B1(n4794), .B2(
        reg_file[689]), .ZN(n6188) );
  AOI22_X1 U5237 ( .A1(n3355), .A2(reg_file[657]), .B1(n4813), .B2(
        reg_file[753]), .ZN(n6189) );
  NAND2_X1 U5238 ( .A1(n6185), .A2(n6373), .ZN(n6204) );
  NAND4_X1 U5239 ( .A1(n6184), .A2(n6183), .A3(n6182), .A4(n6181), .ZN(n6185)
         );
  AOI22_X1 U5240 ( .A1(n3316), .A2(reg_file[17]), .B1(n3315), .B2(reg_file[49]), .ZN(n6181) );
  AOI22_X1 U5241 ( .A1(n3286), .A2(reg_file[113]), .B1(n4805), .B2(
        reg_file[81]), .ZN(n6182) );
  AOI22_X1 U5242 ( .A1(n3314), .A2(reg_file[209]), .B1(n4794), .B2(
        reg_file[177]), .ZN(n6183) );
  AOI22_X1 U5243 ( .A1(n3355), .A2(reg_file[145]), .B1(n4815), .B2(
        reg_file[241]), .ZN(n6184) );
  NAND4_X1 U5244 ( .A1(n5515), .A2(n5514), .A3(n5513), .A4(n5512), .ZN(
        rs2_val_gpr_w[17]) );
  NAND2_X1 U5245 ( .A1(n5511), .A2(n3390), .ZN(n5512) );
  NAND4_X1 U5246 ( .A1(n5510), .A2(n5509), .A3(n5508), .A4(n5507), .ZN(n5511)
         );
  AOI22_X1 U5247 ( .A1(n4788), .A2(reg_file[529]), .B1(n4786), .B2(
        reg_file[561]), .ZN(n5507) );
  AOI22_X1 U5248 ( .A1(n4782), .A2(reg_file[625]), .B1(n4774), .B2(
        reg_file[593]), .ZN(n5508) );
  AOI22_X1 U5249 ( .A1(n3294), .A2(reg_file[689]), .B1(n4765), .B2(
        reg_file[657]), .ZN(n5509) );
  AOI22_X1 U5250 ( .A1(n4756), .A2(reg_file[721]), .B1(n4758), .B2(
        reg_file[753]), .ZN(n5510) );
  NAND2_X1 U5251 ( .A1(n5506), .A2(n3389), .ZN(n5513) );
  NAND4_X1 U5252 ( .A1(n5505), .A2(n5504), .A3(n5503), .A4(n5502), .ZN(n5506)
         );
  AOI22_X1 U5253 ( .A1(n4788), .A2(reg_file[273]), .B1(n4787), .B2(
        reg_file[305]), .ZN(n5502) );
  AOI22_X1 U5254 ( .A1(n4782), .A2(reg_file[369]), .B1(n4774), .B2(
        reg_file[337]), .ZN(n5503) );
  AOI22_X1 U5255 ( .A1(n3294), .A2(reg_file[433]), .B1(n4765), .B2(
        reg_file[401]), .ZN(n5504) );
  AOI22_X1 U5256 ( .A1(n4757), .A2(reg_file[465]), .B1(n4758), .B2(
        reg_file[497]), .ZN(n5505) );
  NAND2_X1 U5257 ( .A1(n5501), .A2(n3361), .ZN(n5514) );
  NAND4_X1 U5258 ( .A1(n5500), .A2(n5499), .A3(n5498), .A4(n5497), .ZN(n5501)
         );
  AOI22_X1 U5259 ( .A1(n4788), .A2(reg_file[785]), .B1(n4787), .B2(
        reg_file[817]), .ZN(n5497) );
  AOI22_X1 U5260 ( .A1(n4782), .A2(reg_file[881]), .B1(n4774), .B2(
        reg_file[849]), .ZN(n5498) );
  AOI22_X1 U5261 ( .A1(n3294), .A2(reg_file[945]), .B1(n4765), .B2(
        reg_file[913]), .ZN(n5499) );
  AOI22_X1 U5262 ( .A1(n4756), .A2(reg_file[977]), .B1(n4758), .B2(
        reg_file[1009]), .ZN(n5500) );
  NAND2_X1 U5263 ( .A1(n5496), .A2(n4754), .ZN(n5515) );
  NAND4_X1 U5264 ( .A1(n5495), .A2(n5494), .A3(n5493), .A4(n5492), .ZN(n5496)
         );
  AOI22_X1 U5265 ( .A1(n4788), .A2(reg_file[17]), .B1(n4787), .B2(reg_file[49]), .ZN(n5492) );
  AOI22_X1 U5266 ( .A1(n4782), .A2(reg_file[113]), .B1(n4774), .B2(
        reg_file[81]), .ZN(n5493) );
  AOI22_X1 U5267 ( .A1(n3294), .A2(reg_file[177]), .B1(n4765), .B2(
        reg_file[145]), .ZN(n5494) );
  AOI22_X1 U5268 ( .A1(n4756), .A2(reg_file[209]), .B1(n4758), .B2(
        reg_file[241]), .ZN(n5495) );
  NAND4_X1 U5269 ( .A1(n6180), .A2(n6179), .A3(n6178), .A4(n6177), .ZN(
        rs1_val_gpr_w[16]) );
  NAND2_X1 U5270 ( .A1(n6176), .A2(n3362), .ZN(n6177) );
  NAND4_X1 U5271 ( .A1(n6175), .A2(n6174), .A3(n6173), .A4(n6172), .ZN(n6176)
         );
  AOI22_X1 U5272 ( .A1(n3316), .A2(reg_file[784]), .B1(n3315), .B2(
        reg_file[816]), .ZN(n6172) );
  AOI22_X1 U5273 ( .A1(n3286), .A2(reg_file[880]), .B1(n4805), .B2(
        reg_file[848]), .ZN(n6173) );
  AOI22_X1 U5274 ( .A1(n3314), .A2(reg_file[976]), .B1(n4794), .B2(
        reg_file[944]), .ZN(n6174) );
  AOI22_X1 U5275 ( .A1(n3386), .A2(reg_file[912]), .B1(n4813), .B2(
        reg_file[1008]), .ZN(n6175) );
  NAND2_X1 U5276 ( .A1(n6171), .A2(n6373), .ZN(n6178) );
  NAND4_X1 U5277 ( .A1(n6170), .A2(n6169), .A3(n6168), .A4(n6167), .ZN(n6171)
         );
  AOI22_X1 U5278 ( .A1(n3316), .A2(reg_file[16]), .B1(n3315), .B2(reg_file[48]), .ZN(n6167) );
  AOI22_X1 U5279 ( .A1(n3285), .A2(reg_file[112]), .B1(n4805), .B2(
        reg_file[80]), .ZN(n6168) );
  AOI22_X1 U5280 ( .A1(n3314), .A2(reg_file[208]), .B1(n4794), .B2(
        reg_file[176]), .ZN(n6169) );
  AOI22_X1 U5281 ( .A1(n3355), .A2(reg_file[144]), .B1(n4813), .B2(
        reg_file[240]), .ZN(n6170) );
  NAND2_X1 U5282 ( .A1(n6166), .A2(n3387), .ZN(n6179) );
  NAND4_X1 U5283 ( .A1(n6165), .A2(n6164), .A3(n6163), .A4(n6162), .ZN(n6166)
         );
  AOI22_X1 U5284 ( .A1(n3316), .A2(reg_file[272]), .B1(n3315), .B2(
        reg_file[304]), .ZN(n6162) );
  AOI22_X1 U5285 ( .A1(n3285), .A2(reg_file[368]), .B1(n4806), .B2(
        reg_file[336]), .ZN(n6163) );
  AOI22_X1 U5286 ( .A1(n3314), .A2(reg_file[464]), .B1(n4794), .B2(
        reg_file[432]), .ZN(n6164) );
  AOI22_X1 U5287 ( .A1(n3386), .A2(reg_file[400]), .B1(n4813), .B2(
        reg_file[496]), .ZN(n6165) );
  NAND2_X1 U5288 ( .A1(n6161), .A2(n3388), .ZN(n6180) );
  NAND4_X1 U5289 ( .A1(n6160), .A2(n6159), .A3(n6158), .A4(n6157), .ZN(n6161)
         );
  AOI22_X1 U5290 ( .A1(n3316), .A2(reg_file[528]), .B1(n3315), .B2(
        reg_file[560]), .ZN(n6157) );
  AOI22_X1 U5291 ( .A1(n3286), .A2(reg_file[624]), .B1(n4805), .B2(
        reg_file[592]), .ZN(n6158) );
  AOI22_X1 U5292 ( .A1(n3314), .A2(reg_file[720]), .B1(n4794), .B2(
        reg_file[688]), .ZN(n6159) );
  AOI22_X1 U5293 ( .A1(n3355), .A2(reg_file[656]), .B1(n4813), .B2(
        reg_file[752]), .ZN(n6160) );
  NAND4_X1 U5294 ( .A1(n5491), .A2(n5490), .A3(n5489), .A4(n5488), .ZN(
        rs2_val_gpr_w[16]) );
  NAND2_X1 U5295 ( .A1(n5487), .A2(n4754), .ZN(n5488) );
  NAND4_X1 U5296 ( .A1(n5486), .A2(n5485), .A3(n5484), .A4(n5483), .ZN(n5487)
         );
  AOI22_X1 U5297 ( .A1(n4788), .A2(reg_file[16]), .B1(n4787), .B2(reg_file[48]), .ZN(n5483) );
  AOI22_X1 U5298 ( .A1(n4782), .A2(reg_file[112]), .B1(n4774), .B2(
        reg_file[80]), .ZN(n5484) );
  AOI22_X1 U5299 ( .A1(n3294), .A2(reg_file[176]), .B1(n4765), .B2(
        reg_file[144]), .ZN(n5485) );
  AOI22_X1 U5300 ( .A1(n4756), .A2(reg_file[208]), .B1(n4758), .B2(
        reg_file[240]), .ZN(n5486) );
  NAND2_X1 U5301 ( .A1(n5482), .A2(n3389), .ZN(n5489) );
  NAND4_X1 U5302 ( .A1(n5481), .A2(n5480), .A3(n5479), .A4(n5478), .ZN(n5482)
         );
  AOI22_X1 U5303 ( .A1(n4788), .A2(reg_file[272]), .B1(n4786), .B2(
        reg_file[304]), .ZN(n5478) );
  AOI22_X1 U5304 ( .A1(n4782), .A2(reg_file[368]), .B1(n4774), .B2(
        reg_file[336]), .ZN(n5479) );
  AOI22_X1 U5305 ( .A1(n3294), .A2(reg_file[432]), .B1(n4765), .B2(
        reg_file[400]), .ZN(n5480) );
  AOI22_X1 U5306 ( .A1(n4757), .A2(reg_file[464]), .B1(n4758), .B2(
        reg_file[496]), .ZN(n5481) );
  NAND2_X1 U5307 ( .A1(n5477), .A2(n3361), .ZN(n5490) );
  NAND4_X1 U5308 ( .A1(n5476), .A2(n5475), .A3(n5474), .A4(n5473), .ZN(n5477)
         );
  AOI22_X1 U5309 ( .A1(n4788), .A2(reg_file[784]), .B1(n4787), .B2(
        reg_file[816]), .ZN(n5473) );
  AOI22_X1 U5310 ( .A1(n4782), .A2(reg_file[880]), .B1(n4774), .B2(
        reg_file[848]), .ZN(n5474) );
  AOI22_X1 U5311 ( .A1(n3294), .A2(reg_file[944]), .B1(n4765), .B2(
        reg_file[912]), .ZN(n5475) );
  AOI22_X1 U5312 ( .A1(n4757), .A2(reg_file[976]), .B1(n4758), .B2(
        reg_file[1008]), .ZN(n5476) );
  NAND2_X1 U5313 ( .A1(n5472), .A2(n3390), .ZN(n5491) );
  NAND4_X1 U5314 ( .A1(n5471), .A2(n5470), .A3(n5469), .A4(n5468), .ZN(n5472)
         );
  AOI22_X1 U5315 ( .A1(n4788), .A2(reg_file[528]), .B1(n4787), .B2(
        reg_file[560]), .ZN(n5468) );
  AOI22_X1 U5316 ( .A1(n4782), .A2(reg_file[624]), .B1(n4774), .B2(
        reg_file[592]), .ZN(n5469) );
  AOI22_X1 U5317 ( .A1(n3294), .A2(reg_file[688]), .B1(n4765), .B2(
        reg_file[656]), .ZN(n5470) );
  AOI22_X1 U5318 ( .A1(n4757), .A2(reg_file[720]), .B1(n4758), .B2(
        reg_file[752]), .ZN(n5471) );
  NAND4_X1 U5319 ( .A1(n6146), .A2(n6145), .A3(n6144), .A4(n6143), .ZN(
        rs1_val_gpr_w[14]) );
  NAND2_X1 U5320 ( .A1(n6142), .A2(n3362), .ZN(n6143) );
  NAND4_X1 U5321 ( .A1(n6141), .A2(n6140), .A3(n6139), .A4(n6138), .ZN(n6142)
         );
  AOI22_X1 U5322 ( .A1(n3316), .A2(reg_file[782]), .B1(n3315), .B2(
        reg_file[814]), .ZN(n6138) );
  AOI22_X1 U5323 ( .A1(n3286), .A2(reg_file[878]), .B1(n3295), .B2(
        reg_file[846]), .ZN(n6139) );
  AOI22_X1 U5324 ( .A1(n3314), .A2(reg_file[974]), .B1(n4793), .B2(
        reg_file[942]), .ZN(n6140) );
  AOI22_X1 U5325 ( .A1(n3355), .A2(reg_file[910]), .B1(n6396), .B2(
        reg_file[1006]), .ZN(n6141) );
  NAND2_X1 U5326 ( .A1(n6137), .A2(n3388), .ZN(n6144) );
  NAND4_X1 U5327 ( .A1(n6136), .A2(n6135), .A3(n6134), .A4(n6133), .ZN(n6137)
         );
  AOI22_X1 U5328 ( .A1(n3316), .A2(reg_file[526]), .B1(n3315), .B2(
        reg_file[558]), .ZN(n6133) );
  AOI22_X1 U5329 ( .A1(n3286), .A2(reg_file[622]), .B1(n3295), .B2(
        reg_file[590]), .ZN(n6134) );
  AOI22_X1 U5330 ( .A1(n3314), .A2(reg_file[718]), .B1(n4793), .B2(
        reg_file[686]), .ZN(n6135) );
  AOI22_X1 U5331 ( .A1(n4790), .A2(reg_file[654]), .B1(n6396), .B2(
        reg_file[750]), .ZN(n6136) );
  NAND2_X1 U5332 ( .A1(n6132), .A2(n3387), .ZN(n6145) );
  NAND4_X1 U5333 ( .A1(n6131), .A2(n6130), .A3(n6129), .A4(n6128), .ZN(n6132)
         );
  AOI22_X1 U5334 ( .A1(n3316), .A2(reg_file[270]), .B1(n3315), .B2(
        reg_file[302]), .ZN(n6128) );
  AOI22_X1 U5335 ( .A1(n3285), .A2(reg_file[366]), .B1(n3295), .B2(
        reg_file[334]), .ZN(n6129) );
  AOI22_X1 U5336 ( .A1(n3314), .A2(reg_file[462]), .B1(n4793), .B2(
        reg_file[430]), .ZN(n6130) );
  AOI22_X1 U5337 ( .A1(n3355), .A2(reg_file[398]), .B1(n6396), .B2(
        reg_file[494]), .ZN(n6131) );
  NAND2_X1 U5338 ( .A1(n6127), .A2(n6373), .ZN(n6146) );
  NAND4_X1 U5339 ( .A1(n6126), .A2(n6125), .A3(n6124), .A4(n6123), .ZN(n6127)
         );
  AOI22_X1 U5340 ( .A1(n3316), .A2(reg_file[14]), .B1(n3315), .B2(reg_file[46]), .ZN(n6123) );
  AOI22_X1 U5341 ( .A1(n3285), .A2(reg_file[110]), .B1(n3295), .B2(
        reg_file[78]), .ZN(n6124) );
  AOI22_X1 U5342 ( .A1(n3314), .A2(reg_file[206]), .B1(n4793), .B2(
        reg_file[174]), .ZN(n6125) );
  AOI22_X1 U5343 ( .A1(n3386), .A2(reg_file[142]), .B1(n6396), .B2(
        reg_file[238]), .ZN(n6126) );
  NAND4_X1 U5344 ( .A1(n5454), .A2(n5453), .A3(n5452), .A4(n5451), .ZN(n5455)
         );
  AOI22_X1 U5345 ( .A1(n4789), .A2(reg_file[526]), .B1(n4787), .B2(
        reg_file[558]), .ZN(n5451) );
  AOI22_X1 U5346 ( .A1(n4783), .A2(reg_file[622]), .B1(n4773), .B2(
        reg_file[590]), .ZN(n5452) );
  AOI22_X1 U5347 ( .A1(n3294), .A2(reg_file[686]), .B1(n4764), .B2(
        reg_file[654]), .ZN(n5453) );
  AOI22_X1 U5348 ( .A1(n4757), .A2(reg_file[718]), .B1(n4758), .B2(
        reg_file[750]), .ZN(n5454) );
  AOI22_X1 U5349 ( .A1(n4789), .A2(reg_file[270]), .B1(n4787), .B2(
        reg_file[302]), .ZN(n5447) );
  AOI22_X1 U5350 ( .A1(n4784), .A2(reg_file[366]), .B1(n4773), .B2(
        reg_file[334]), .ZN(n5448) );
  AOI22_X1 U5351 ( .A1(n3294), .A2(reg_file[430]), .B1(n4764), .B2(
        reg_file[398]), .ZN(n5449) );
  AOI22_X1 U5352 ( .A1(n4755), .A2(reg_file[462]), .B1(n4758), .B2(
        reg_file[494]), .ZN(n5450) );
  AOI22_X1 U5353 ( .A1(n4789), .A2(reg_file[782]), .B1(n4786), .B2(
        reg_file[814]), .ZN(n5443) );
  AOI22_X1 U5354 ( .A1(n4783), .A2(reg_file[878]), .B1(n4773), .B2(
        reg_file[846]), .ZN(n5444) );
  AOI22_X1 U5355 ( .A1(n3294), .A2(reg_file[942]), .B1(n4764), .B2(
        reg_file[910]), .ZN(n5445) );
  AOI22_X1 U5356 ( .A1(n4757), .A2(reg_file[974]), .B1(n4758), .B2(
        reg_file[1006]), .ZN(n5446) );
  AOI22_X1 U5357 ( .A1(n3296), .A2(reg_file[14]), .B1(n4787), .B2(reg_file[46]), .ZN(n5439) );
  AOI22_X1 U5358 ( .A1(n5811), .A2(reg_file[110]), .B1(n4773), .B2(
        reg_file[78]), .ZN(n5440) );
  AOI22_X1 U5359 ( .A1(n3294), .A2(reg_file[174]), .B1(n4764), .B2(
        reg_file[142]), .ZN(n5441) );
  AOI22_X1 U5360 ( .A1(n4755), .A2(reg_file[206]), .B1(n4758), .B2(
        reg_file[238]), .ZN(n5442) );
  NAND2_X1 U5361 ( .A1(n6118), .A2(n3362), .ZN(n6119) );
  NAND4_X1 U5362 ( .A1(n6117), .A2(n6116), .A3(n6115), .A4(n6114), .ZN(n6118)
         );
  AOI22_X1 U5363 ( .A1(n3316), .A2(reg_file[781]), .B1(n3315), .B2(
        reg_file[813]), .ZN(n6114) );
  AOI22_X1 U5364 ( .A1(n3286), .A2(reg_file[877]), .B1(n3295), .B2(
        reg_file[845]), .ZN(n6115) );
  AOI22_X1 U5365 ( .A1(n3314), .A2(reg_file[973]), .B1(n4793), .B2(
        reg_file[941]), .ZN(n6116) );
  AOI22_X1 U5366 ( .A1(n3355), .A2(reg_file[909]), .B1(n4815), .B2(
        reg_file[1005]), .ZN(n6117) );
  NAND2_X1 U5367 ( .A1(n6113), .A2(n3387), .ZN(n6120) );
  NAND4_X1 U5368 ( .A1(n6112), .A2(n6111), .A3(n6110), .A4(n6109), .ZN(n6113)
         );
  AOI22_X1 U5369 ( .A1(n3316), .A2(reg_file[269]), .B1(n3315), .B2(
        reg_file[301]), .ZN(n6109) );
  AOI22_X1 U5370 ( .A1(n3286), .A2(reg_file[365]), .B1(n3295), .B2(
        reg_file[333]), .ZN(n6110) );
  AOI22_X1 U5371 ( .A1(n3314), .A2(reg_file[461]), .B1(n4793), .B2(
        reg_file[429]), .ZN(n6111) );
  AOI22_X1 U5372 ( .A1(n3355), .A2(reg_file[397]), .B1(n4815), .B2(
        reg_file[493]), .ZN(n6112) );
  NAND2_X1 U5373 ( .A1(n6108), .A2(n3388), .ZN(n6121) );
  NAND4_X1 U5374 ( .A1(n6107), .A2(n6106), .A3(n6105), .A4(n6104), .ZN(n6108)
         );
  AOI22_X1 U5375 ( .A1(n3316), .A2(reg_file[525]), .B1(n3315), .B2(
        reg_file[557]), .ZN(n6104) );
  AOI22_X1 U5376 ( .A1(n3285), .A2(reg_file[621]), .B1(n3295), .B2(
        reg_file[589]), .ZN(n6105) );
  AOI22_X1 U5377 ( .A1(n3314), .A2(reg_file[717]), .B1(n4793), .B2(
        reg_file[685]), .ZN(n6106) );
  AOI22_X1 U5378 ( .A1(n3355), .A2(reg_file[653]), .B1(n6396), .B2(
        reg_file[749]), .ZN(n6107) );
  NAND2_X1 U5379 ( .A1(n6103), .A2(n6373), .ZN(n6122) );
  NAND4_X1 U5380 ( .A1(n6102), .A2(n6101), .A3(n6100), .A4(n6099), .ZN(n6103)
         );
  AOI22_X1 U5381 ( .A1(n3316), .A2(reg_file[13]), .B1(n3315), .B2(reg_file[45]), .ZN(n6099) );
  AOI22_X1 U5382 ( .A1(n3286), .A2(reg_file[109]), .B1(n3295), .B2(
        reg_file[77]), .ZN(n6100) );
  AOI22_X1 U5383 ( .A1(n3314), .A2(reg_file[205]), .B1(n4793), .B2(
        reg_file[173]), .ZN(n6101) );
  AOI22_X1 U5384 ( .A1(n3355), .A2(reg_file[141]), .B1(n6396), .B2(
        reg_file[237]), .ZN(n6102) );
  AOI22_X1 U5385 ( .A1(n4789), .A2(reg_file[525]), .B1(n4787), .B2(
        reg_file[557]), .ZN(n5435) );
  AOI22_X1 U5386 ( .A1(n4783), .A2(reg_file[621]), .B1(n4773), .B2(
        reg_file[589]), .ZN(n5436) );
  AOI22_X1 U5387 ( .A1(n3294), .A2(reg_file[685]), .B1(n4764), .B2(
        reg_file[653]), .ZN(n5437) );
  AOI22_X1 U5388 ( .A1(n4756), .A2(reg_file[717]), .B1(n4758), .B2(
        reg_file[749]), .ZN(n5438) );
  AOI22_X1 U5389 ( .A1(n4789), .A2(reg_file[269]), .B1(n4786), .B2(
        reg_file[301]), .ZN(n5431) );
  AOI22_X1 U5390 ( .A1(n4783), .A2(reg_file[365]), .B1(n4773), .B2(
        reg_file[333]), .ZN(n5432) );
  AOI22_X1 U5391 ( .A1(n3294), .A2(reg_file[429]), .B1(n4764), .B2(
        reg_file[397]), .ZN(n5433) );
  AOI22_X1 U5392 ( .A1(n4755), .A2(reg_file[461]), .B1(n4758), .B2(
        reg_file[493]), .ZN(n5434) );
  AOI22_X1 U5393 ( .A1(n4789), .A2(reg_file[781]), .B1(n4786), .B2(
        reg_file[813]), .ZN(n5427) );
  AOI22_X1 U5394 ( .A1(n4783), .A2(reg_file[877]), .B1(n4773), .B2(
        reg_file[845]), .ZN(n5428) );
  AOI22_X1 U5395 ( .A1(n3294), .A2(reg_file[941]), .B1(n4764), .B2(
        reg_file[909]), .ZN(n5429) );
  AOI22_X1 U5396 ( .A1(n4757), .A2(reg_file[973]), .B1(n4758), .B2(
        reg_file[1005]), .ZN(n5430) );
  AOI22_X1 U5397 ( .A1(n4789), .A2(reg_file[13]), .B1(n4786), .B2(reg_file[45]), .ZN(n5425) );
  AOI22_X1 U5398 ( .A1(n4757), .A2(reg_file[205]), .B1(n4758), .B2(
        reg_file[237]), .ZN(n5426) );
  NAND2_X1 U5399 ( .A1(n6094), .A2(n3362), .ZN(n6095) );
  NAND4_X1 U5400 ( .A1(n6093), .A2(n6092), .A3(n6091), .A4(n6090), .ZN(n6094)
         );
  AOI22_X1 U5401 ( .A1(n3316), .A2(reg_file[780]), .B1(n3315), .B2(
        reg_file[812]), .ZN(n6090) );
  AOI22_X1 U5402 ( .A1(n3285), .A2(reg_file[876]), .B1(n3295), .B2(
        reg_file[844]), .ZN(n6091) );
  AOI22_X1 U5403 ( .A1(n3314), .A2(reg_file[972]), .B1(n4793), .B2(
        reg_file[940]), .ZN(n6092) );
  AOI22_X1 U5404 ( .A1(reg_file[908]), .A2(n3386), .B1(n4815), .B2(
        reg_file[1004]), .ZN(n6093) );
  NAND2_X1 U5405 ( .A1(n6089), .A2(n3388), .ZN(n6096) );
  NAND4_X1 U5406 ( .A1(n6088), .A2(n6087), .A3(n6086), .A4(n6085), .ZN(n6089)
         );
  AOI22_X1 U5407 ( .A1(n3316), .A2(reg_file[524]), .B1(n3315), .B2(
        reg_file[556]), .ZN(n6085) );
  AOI22_X1 U5408 ( .A1(n3285), .A2(reg_file[620]), .B1(n3295), .B2(
        reg_file[588]), .ZN(n6086) );
  AOI22_X1 U5409 ( .A1(n3314), .A2(reg_file[716]), .B1(n4793), .B2(
        reg_file[684]), .ZN(n6087) );
  AOI22_X1 U5410 ( .A1(reg_file[652]), .A2(n3386), .B1(n4815), .B2(
        reg_file[748]), .ZN(n6088) );
  NAND2_X1 U5411 ( .A1(n6084), .A2(n3387), .ZN(n6097) );
  NAND4_X1 U5412 ( .A1(n6083), .A2(n6082), .A3(n6081), .A4(n6080), .ZN(n6084)
         );
  AOI22_X1 U5413 ( .A1(n3316), .A2(reg_file[268]), .B1(n3315), .B2(
        reg_file[300]), .ZN(n6080) );
  AOI22_X1 U5414 ( .A1(n3285), .A2(reg_file[364]), .B1(n3295), .B2(
        reg_file[332]), .ZN(n6081) );
  AOI22_X1 U5415 ( .A1(n3314), .A2(reg_file[460]), .B1(n4793), .B2(
        reg_file[428]), .ZN(n6082) );
  AOI22_X1 U5416 ( .A1(n3386), .A2(reg_file[396]), .B1(n4815), .B2(
        reg_file[492]), .ZN(n6083) );
  NAND2_X1 U5417 ( .A1(n6079), .A2(n6373), .ZN(n6098) );
  NAND4_X1 U5418 ( .A1(n6078), .A2(n6077), .A3(n6076), .A4(n6075), .ZN(n6079)
         );
  AOI22_X1 U5419 ( .A1(n3316), .A2(reg_file[12]), .B1(n3315), .B2(reg_file[44]), .ZN(n6075) );
  AOI22_X1 U5420 ( .A1(n3286), .A2(reg_file[108]), .B1(n3295), .B2(
        reg_file[76]), .ZN(n6076) );
  AOI22_X1 U5421 ( .A1(n3314), .A2(reg_file[204]), .B1(n4793), .B2(
        reg_file[172]), .ZN(n6077) );
  AOI22_X1 U5422 ( .A1(reg_file[140]), .A2(n3355), .B1(n4815), .B2(
        reg_file[236]), .ZN(n6078) );
  NAND4_X1 U5423 ( .A1(n5423), .A2(n5422), .A3(n5421), .A4(n5420), .ZN(n5424)
         );
  AOI22_X1 U5424 ( .A1(n4789), .A2(reg_file[780]), .B1(n4787), .B2(
        reg_file[812]), .ZN(n5420) );
  AOI22_X1 U5425 ( .A1(n4783), .A2(reg_file[876]), .B1(n4773), .B2(
        reg_file[844]), .ZN(n5421) );
  AOI22_X1 U5426 ( .A1(n3294), .A2(reg_file[940]), .B1(n4764), .B2(
        reg_file[908]), .ZN(n5422) );
  AOI22_X1 U5427 ( .A1(n4757), .A2(reg_file[972]), .B1(n4759), .B2(
        reg_file[1004]), .ZN(n5423) );
  NAND4_X1 U5428 ( .A1(n5418), .A2(n5417), .A3(n5416), .A4(n5415), .ZN(n5419)
         );
  AOI22_X1 U5429 ( .A1(n4789), .A2(reg_file[524]), .B1(n4786), .B2(
        reg_file[556]), .ZN(n5415) );
  AOI22_X1 U5430 ( .A1(n4784), .A2(reg_file[620]), .B1(n4773), .B2(
        reg_file[588]), .ZN(n5416) );
  AOI22_X1 U5431 ( .A1(n3294), .A2(reg_file[684]), .B1(n4764), .B2(
        reg_file[652]), .ZN(n5417) );
  AOI22_X1 U5432 ( .A1(n4755), .A2(reg_file[716]), .B1(n4759), .B2(
        reg_file[748]), .ZN(n5418) );
  AOI22_X1 U5433 ( .A1(n4789), .A2(reg_file[12]), .B1(n4786), .B2(reg_file[44]), .ZN(n5411) );
  AOI22_X1 U5434 ( .A1(n4783), .A2(reg_file[108]), .B1(n4773), .B2(
        reg_file[76]), .ZN(n5412) );
  AOI22_X1 U5435 ( .A1(n3294), .A2(reg_file[172]), .B1(n4764), .B2(
        reg_file[140]), .ZN(n5413) );
  AOI22_X1 U5436 ( .A1(n4757), .A2(reg_file[204]), .B1(n4759), .B2(
        reg_file[236]), .ZN(n5414) );
  AOI22_X1 U5437 ( .A1(n4789), .A2(reg_file[268]), .B1(n4786), .B2(
        reg_file[300]), .ZN(n5407) );
  AOI22_X1 U5438 ( .A1(n4783), .A2(reg_file[364]), .B1(n4773), .B2(
        reg_file[332]), .ZN(n5408) );
  AOI22_X1 U5439 ( .A1(n3294), .A2(reg_file[428]), .B1(n4764), .B2(
        reg_file[396]), .ZN(n5409) );
  AOI22_X1 U5440 ( .A1(n4757), .A2(reg_file[460]), .B1(n4759), .B2(
        reg_file[492]), .ZN(n5410) );
  NAND2_X1 U5441 ( .A1(n6070), .A2(n3362), .ZN(n6071) );
  NAND4_X1 U5442 ( .A1(n6069), .A2(n6068), .A3(n6067), .A4(n6066), .ZN(n6070)
         );
  AOI22_X1 U5443 ( .A1(n4812), .A2(reg_file[779]), .B1(n4808), .B2(
        reg_file[811]), .ZN(n6066) );
  AOI22_X1 U5444 ( .A1(n3285), .A2(reg_file[875]), .B1(n3295), .B2(
        reg_file[843]), .ZN(n6067) );
  AOI22_X1 U5445 ( .A1(n4799), .A2(reg_file[971]), .B1(n4792), .B2(
        reg_file[939]), .ZN(n6068) );
  AOI22_X1 U5446 ( .A1(n3355), .A2(reg_file[907]), .B1(n4815), .B2(
        reg_file[1003]), .ZN(n6069) );
  NAND2_X1 U5447 ( .A1(n6065), .A2(n6392), .ZN(n6072) );
  NAND4_X1 U5448 ( .A1(n6064), .A2(n6063), .A3(n6062), .A4(n6061), .ZN(n6065)
         );
  AOI22_X1 U5449 ( .A1(n4812), .A2(reg_file[523]), .B1(n4808), .B2(
        reg_file[555]), .ZN(n6061) );
  AOI22_X1 U5450 ( .A1(n3285), .A2(reg_file[619]), .B1(n3295), .B2(
        reg_file[587]), .ZN(n6062) );
  AOI22_X1 U5451 ( .A1(n4799), .A2(reg_file[715]), .B1(n4792), .B2(
        reg_file[683]), .ZN(n6063) );
  AOI22_X1 U5452 ( .A1(n4790), .A2(reg_file[651]), .B1(n4815), .B2(
        reg_file[747]), .ZN(n6064) );
  NAND2_X1 U5453 ( .A1(n6060), .A2(n6381), .ZN(n6073) );
  NAND4_X1 U5454 ( .A1(n6059), .A2(n6058), .A3(n6057), .A4(n6056), .ZN(n6060)
         );
  AOI22_X1 U5455 ( .A1(n4812), .A2(reg_file[267]), .B1(n4808), .B2(
        reg_file[299]), .ZN(n6056) );
  AOI22_X1 U5456 ( .A1(n3285), .A2(reg_file[363]), .B1(n3295), .B2(
        reg_file[331]), .ZN(n6057) );
  AOI22_X1 U5457 ( .A1(n4799), .A2(reg_file[459]), .B1(n4792), .B2(
        reg_file[427]), .ZN(n6058) );
  AOI22_X1 U5458 ( .A1(n3386), .A2(reg_file[395]), .B1(n4815), .B2(
        reg_file[491]), .ZN(n6059) );
  NAND2_X1 U5459 ( .A1(n6055), .A2(n6373), .ZN(n6074) );
  NAND4_X1 U5460 ( .A1(n6054), .A2(n6053), .A3(n6052), .A4(n6051), .ZN(n6055)
         );
  AOI22_X1 U5461 ( .A1(n4812), .A2(reg_file[11]), .B1(n4808), .B2(reg_file[43]), .ZN(n6051) );
  AOI22_X1 U5462 ( .A1(n3286), .A2(reg_file[107]), .B1(n3295), .B2(
        reg_file[75]), .ZN(n6052) );
  AOI22_X1 U5463 ( .A1(n4799), .A2(reg_file[203]), .B1(n4792), .B2(
        reg_file[171]), .ZN(n6053) );
  AOI22_X1 U5464 ( .A1(n4790), .A2(reg_file[139]), .B1(n4815), .B2(
        reg_file[235]), .ZN(n6054) );
  NAND2_X1 U5465 ( .A1(n5402), .A2(n3361), .ZN(n5403) );
  NAND4_X1 U5466 ( .A1(n5401), .A2(n5400), .A3(n5399), .A4(n5398), .ZN(n5402)
         );
  AOI22_X1 U5467 ( .A1(n4789), .A2(reg_file[779]), .B1(n4786), .B2(
        reg_file[811]), .ZN(n5398) );
  AOI22_X1 U5468 ( .A1(n4783), .A2(reg_file[875]), .B1(n4772), .B2(
        reg_file[843]), .ZN(n5399) );
  AOI22_X1 U5469 ( .A1(n3294), .A2(reg_file[939]), .B1(n3769), .B2(
        reg_file[907]), .ZN(n5400) );
  AOI22_X1 U5470 ( .A1(n4756), .A2(reg_file[971]), .B1(n4759), .B2(
        reg_file[1003]), .ZN(n5401) );
  NAND2_X1 U5471 ( .A1(n5397), .A2(n3389), .ZN(n5404) );
  NAND4_X1 U5472 ( .A1(n5396), .A2(n5395), .A3(n5394), .A4(n5393), .ZN(n5397)
         );
  AOI22_X1 U5473 ( .A1(n4789), .A2(reg_file[267]), .B1(n4786), .B2(
        reg_file[299]), .ZN(n5393) );
  AOI22_X1 U5474 ( .A1(n4783), .A2(reg_file[363]), .B1(n4772), .B2(
        reg_file[331]), .ZN(n5394) );
  AOI22_X1 U5475 ( .A1(n3294), .A2(reg_file[427]), .B1(n4766), .B2(
        reg_file[395]), .ZN(n5395) );
  AOI22_X1 U5476 ( .A1(n4756), .A2(reg_file[459]), .B1(n4759), .B2(
        reg_file[491]), .ZN(n5396) );
  NAND2_X1 U5477 ( .A1(n5392), .A2(n3390), .ZN(n5405) );
  NAND4_X1 U5478 ( .A1(n5391), .A2(n5390), .A3(n5389), .A4(n5388), .ZN(n5392)
         );
  AOI22_X1 U5479 ( .A1(n4789), .A2(reg_file[523]), .B1(n4786), .B2(
        reg_file[555]), .ZN(n5388) );
  AOI22_X1 U5480 ( .A1(n4783), .A2(reg_file[619]), .B1(n4772), .B2(
        reg_file[587]), .ZN(n5389) );
  AOI22_X1 U5481 ( .A1(n3294), .A2(reg_file[683]), .B1(n4767), .B2(
        reg_file[651]), .ZN(n5390) );
  AOI22_X1 U5482 ( .A1(n4757), .A2(reg_file[715]), .B1(n4759), .B2(
        reg_file[747]), .ZN(n5391) );
  NAND2_X1 U5483 ( .A1(n5387), .A2(n5805), .ZN(n5406) );
  NAND4_X1 U5484 ( .A1(n5386), .A2(n5385), .A3(n5384), .A4(n5383), .ZN(n5387)
         );
  AOI22_X1 U5485 ( .A1(n4789), .A2(reg_file[11]), .B1(n4786), .B2(reg_file[43]), .ZN(n5383) );
  AOI22_X1 U5486 ( .A1(n4783), .A2(reg_file[107]), .B1(n4772), .B2(
        reg_file[75]), .ZN(n5384) );
  AOI22_X1 U5487 ( .A1(n3294), .A2(reg_file[171]), .B1(n4768), .B2(
        reg_file[139]), .ZN(n5385) );
  AOI22_X1 U5488 ( .A1(n4757), .A2(reg_file[203]), .B1(n4759), .B2(
        reg_file[235]), .ZN(n5386) );
  NAND2_X1 U5489 ( .A1(n6046), .A2(n6381), .ZN(n6047) );
  NAND4_X1 U5490 ( .A1(n6045), .A2(n6044), .A3(n6043), .A4(n6042), .ZN(n6046)
         );
  AOI22_X1 U5491 ( .A1(n4812), .A2(reg_file[266]), .B1(n4808), .B2(
        reg_file[298]), .ZN(n6042) );
  AOI22_X1 U5492 ( .A1(n3286), .A2(reg_file[362]), .B1(n3295), .B2(
        reg_file[330]), .ZN(n6043) );
  AOI22_X1 U5493 ( .A1(n4799), .A2(reg_file[458]), .B1(n4792), .B2(
        reg_file[426]), .ZN(n6044) );
  AOI22_X1 U5494 ( .A1(n4790), .A2(reg_file[394]), .B1(n4815), .B2(
        reg_file[490]), .ZN(n6045) );
  NAND2_X1 U5495 ( .A1(n6041), .A2(n6392), .ZN(n6048) );
  NAND4_X1 U5496 ( .A1(n6040), .A2(n6039), .A3(n6038), .A4(n6037), .ZN(n6041)
         );
  AOI22_X1 U5497 ( .A1(n4812), .A2(reg_file[522]), .B1(n4808), .B2(
        reg_file[554]), .ZN(n6037) );
  AOI22_X1 U5498 ( .A1(n3286), .A2(reg_file[618]), .B1(n3295), .B2(
        reg_file[586]), .ZN(n6038) );
  AOI22_X1 U5499 ( .A1(n4799), .A2(reg_file[714]), .B1(n4792), .B2(
        reg_file[682]), .ZN(n6039) );
  AOI22_X1 U5500 ( .A1(n3355), .A2(reg_file[650]), .B1(n4815), .B2(
        reg_file[746]), .ZN(n6040) );
  NAND2_X1 U5501 ( .A1(n6036), .A2(n3362), .ZN(n6049) );
  NAND4_X1 U5502 ( .A1(n6035), .A2(n6034), .A3(n6033), .A4(n6032), .ZN(n6036)
         );
  AOI22_X1 U5503 ( .A1(n4812), .A2(reg_file[778]), .B1(n4808), .B2(
        reg_file[810]), .ZN(n6032) );
  AOI22_X1 U5504 ( .A1(n3286), .A2(reg_file[874]), .B1(n3295), .B2(
        reg_file[842]), .ZN(n6033) );
  AOI22_X1 U5505 ( .A1(n4799), .A2(reg_file[970]), .B1(n4792), .B2(
        reg_file[938]), .ZN(n6034) );
  AOI22_X1 U5506 ( .A1(n4790), .A2(reg_file[906]), .B1(n4815), .B2(
        reg_file[1002]), .ZN(n6035) );
  NAND2_X1 U5507 ( .A1(n6031), .A2(n6373), .ZN(n6050) );
  NAND4_X1 U5508 ( .A1(n6030), .A2(n6029), .A3(n6028), .A4(n6027), .ZN(n6031)
         );
  AOI22_X1 U5509 ( .A1(n4812), .A2(reg_file[10]), .B1(n4808), .B2(reg_file[42]), .ZN(n6027) );
  AOI22_X1 U5510 ( .A1(n3286), .A2(reg_file[106]), .B1(n3295), .B2(
        reg_file[74]), .ZN(n6028) );
  AOI22_X1 U5511 ( .A1(n4799), .A2(reg_file[202]), .B1(n4792), .B2(
        reg_file[170]), .ZN(n6029) );
  AOI22_X1 U5512 ( .A1(n3355), .A2(reg_file[138]), .B1(n4815), .B2(
        reg_file[234]), .ZN(n6030) );
  NAND4_X1 U5513 ( .A1(n5381), .A2(n5380), .A3(n5379), .A4(n5378), .ZN(n5382)
         );
  AOI22_X1 U5514 ( .A1(n4789), .A2(reg_file[522]), .B1(n4787), .B2(
        reg_file[554]), .ZN(n5378) );
  AOI22_X1 U5515 ( .A1(n4783), .A2(reg_file[618]), .B1(n4772), .B2(
        reg_file[586]), .ZN(n5379) );
  AOI22_X1 U5516 ( .A1(n3294), .A2(reg_file[682]), .B1(n3769), .B2(
        reg_file[650]), .ZN(n5380) );
  AOI22_X1 U5517 ( .A1(n3519), .A2(reg_file[714]), .B1(n4759), .B2(
        reg_file[746]), .ZN(n5381) );
  NAND4_X1 U5518 ( .A1(n5376), .A2(n5375), .A3(n5374), .A4(n5373), .ZN(n5377)
         );
  AOI22_X1 U5519 ( .A1(n4789), .A2(reg_file[266]), .B1(n4787), .B2(
        reg_file[298]), .ZN(n5373) );
  AOI22_X1 U5520 ( .A1(n4783), .A2(reg_file[362]), .B1(n4772), .B2(
        reg_file[330]), .ZN(n5374) );
  AOI22_X1 U5521 ( .A1(n3294), .A2(reg_file[426]), .B1(n3769), .B2(
        reg_file[394]), .ZN(n5375) );
  AOI22_X1 U5522 ( .A1(n4755), .A2(reg_file[458]), .B1(n4759), .B2(
        reg_file[490]), .ZN(n5376) );
  NAND4_X1 U5523 ( .A1(n5371), .A2(n5370), .A3(n5369), .A4(n5368), .ZN(n5372)
         );
  AOI22_X1 U5524 ( .A1(n4789), .A2(reg_file[778]), .B1(n4787), .B2(
        reg_file[810]), .ZN(n5368) );
  AOI22_X1 U5525 ( .A1(n4783), .A2(reg_file[874]), .B1(n4772), .B2(
        reg_file[842]), .ZN(n5369) );
  AOI22_X1 U5526 ( .A1(n3294), .A2(reg_file[938]), .B1(n4766), .B2(
        reg_file[906]), .ZN(n5370) );
  BUF_X1 U5527 ( .A(n3769), .Z(n4766) );
  AOI22_X1 U5528 ( .A1(n4757), .A2(reg_file[970]), .B1(n4759), .B2(
        reg_file[1002]), .ZN(n5371) );
  AOI22_X1 U5529 ( .A1(n4789), .A2(reg_file[10]), .B1(n4786), .B2(reg_file[42]), .ZN(n5364) );
  AOI22_X1 U5530 ( .A1(n4783), .A2(reg_file[106]), .B1(n4772), .B2(
        reg_file[74]), .ZN(n5365) );
  AOI22_X1 U5531 ( .A1(n3294), .A2(reg_file[170]), .B1(n4767), .B2(
        reg_file[138]), .ZN(n5366) );
  AOI22_X1 U5532 ( .A1(n4757), .A2(reg_file[202]), .B1(n4759), .B2(
        reg_file[234]), .ZN(n5367) );
  AOI22_X1 U5533 ( .A1(n3316), .A2(reg_file[271]), .B1(n3315), .B2(
        reg_file[303]), .ZN(n6153) );
  AOI22_X1 U5534 ( .A1(n3286), .A2(reg_file[367]), .B1(n3359), .B2(
        reg_file[335]), .ZN(n6154) );
  AOI22_X1 U5535 ( .A1(n3314), .A2(reg_file[463]), .B1(n4794), .B2(
        reg_file[431]), .ZN(n6155) );
  AOI22_X1 U5536 ( .A1(n4790), .A2(reg_file[399]), .B1(n4815), .B2(
        reg_file[495]), .ZN(n6156) );
  AOI22_X1 U5537 ( .A1(n3316), .A2(reg_file[15]), .B1(n3315), .B2(reg_file[47]), .ZN(n6149) );
  AOI22_X1 U5538 ( .A1(n3286), .A2(reg_file[111]), .B1(n3359), .B2(
        reg_file[79]), .ZN(n6150) );
  AOI22_X1 U5539 ( .A1(n3314), .A2(reg_file[207]), .B1(n4794), .B2(
        reg_file[175]), .ZN(n6151) );
  AOI22_X1 U5540 ( .A1(n3355), .A2(reg_file[143]), .B1(n4815), .B2(
        reg_file[239]), .ZN(n6152) );
  AOI22_X1 U5541 ( .A1(n3314), .A2(reg_file[975]), .B1(n4794), .B2(
        reg_file[943]), .ZN(n6147) );
  AOI22_X1 U5542 ( .A1(n4790), .A2(reg_file[911]), .B1(n4814), .B2(
        reg_file[1007]), .ZN(n6148) );
  AOI22_X1 U5543 ( .A1(n4788), .A2(reg_file[783]), .B1(n4787), .B2(
        reg_file[815]), .ZN(n5464) );
  AOI22_X1 U5544 ( .A1(n4782), .A2(reg_file[879]), .B1(n4774), .B2(
        reg_file[847]), .ZN(n5465) );
  AOI22_X1 U5545 ( .A1(n3294), .A2(reg_file[943]), .B1(n4765), .B2(
        reg_file[911]), .ZN(n5466) );
  AOI22_X1 U5546 ( .A1(n4755), .A2(reg_file[975]), .B1(n4758), .B2(
        reg_file[1007]), .ZN(n5467) );
  AOI22_X1 U5547 ( .A1(n4789), .A2(reg_file[527]), .B1(n4787), .B2(
        reg_file[559]), .ZN(n5460) );
  AOI22_X1 U5548 ( .A1(n4784), .A2(reg_file[623]), .B1(n4774), .B2(
        reg_file[591]), .ZN(n5461) );
  AOI22_X1 U5549 ( .A1(n3294), .A2(reg_file[687]), .B1(n4765), .B2(
        reg_file[655]), .ZN(n5462) );
  AOI22_X1 U5550 ( .A1(n4756), .A2(reg_file[719]), .B1(n4758), .B2(
        reg_file[751]), .ZN(n5463) );
  AOI22_X1 U5551 ( .A1(n3296), .A2(reg_file[15]), .B1(n4786), .B2(reg_file[47]), .ZN(n5456) );
  AOI22_X1 U5552 ( .A1(n4783), .A2(reg_file[111]), .B1(n4774), .B2(
        reg_file[79]), .ZN(n5457) );
  AOI22_X1 U5553 ( .A1(n3294), .A2(reg_file[175]), .B1(n4765), .B2(
        reg_file[143]), .ZN(n5458) );
  AOI22_X1 U5554 ( .A1(n4757), .A2(reg_file[207]), .B1(n4758), .B2(
        reg_file[239]), .ZN(n5459) );
  NAND2_X1 U5555 ( .A1(n5998), .A2(n3362), .ZN(n5999) );
  NAND4_X1 U5556 ( .A1(n5997), .A2(n5996), .A3(n5995), .A4(n5994), .ZN(n5998)
         );
  AOI22_X1 U5557 ( .A1(n3358), .A2(reg_file[776]), .B1(n4809), .B2(
        reg_file[808]), .ZN(n5994) );
  AOI22_X1 U5558 ( .A1(n3286), .A2(reg_file[872]), .B1(n4804), .B2(
        reg_file[840]), .ZN(n5995) );
  AOI22_X1 U5559 ( .A1(n4800), .A2(reg_file[968]), .B1(n4797), .B2(
        reg_file[936]), .ZN(n5996) );
  AOI22_X1 U5560 ( .A1(n4790), .A2(reg_file[904]), .B1(n4815), .B2(
        reg_file[1000]), .ZN(n5997) );
  NAND2_X1 U5561 ( .A1(n5993), .A2(n6373), .ZN(n6000) );
  NAND4_X1 U5562 ( .A1(n5992), .A2(n5991), .A3(n5990), .A4(n5989), .ZN(n5993)
         );
  AOI22_X1 U5563 ( .A1(n3358), .A2(reg_file[8]), .B1(n4809), .B2(reg_file[40]), 
        .ZN(n5989) );
  AOI22_X1 U5564 ( .A1(n3285), .A2(reg_file[104]), .B1(n4804), .B2(
        reg_file[72]), .ZN(n5990) );
  AOI22_X1 U5565 ( .A1(n4799), .A2(reg_file[200]), .B1(n4797), .B2(
        reg_file[168]), .ZN(n5991) );
  AOI22_X1 U5566 ( .A1(n3355), .A2(reg_file[136]), .B1(n4815), .B2(
        reg_file[232]), .ZN(n5992) );
  NAND2_X1 U5567 ( .A1(n5988), .A2(n6381), .ZN(n6001) );
  NAND4_X1 U5568 ( .A1(n5987), .A2(n5986), .A3(n5985), .A4(n5984), .ZN(n5988)
         );
  AOI22_X1 U5569 ( .A1(n4811), .A2(reg_file[264]), .B1(n4809), .B2(
        reg_file[296]), .ZN(n5984) );
  AOI22_X1 U5570 ( .A1(n3285), .A2(reg_file[360]), .B1(n4804), .B2(
        reg_file[328]), .ZN(n5985) );
  AOI22_X1 U5571 ( .A1(n4798), .A2(reg_file[456]), .B1(n4796), .B2(
        reg_file[424]), .ZN(n5986) );
  AOI22_X1 U5572 ( .A1(n3355), .A2(reg_file[392]), .B1(n4815), .B2(
        reg_file[488]), .ZN(n5987) );
  NAND2_X1 U5573 ( .A1(n5983), .A2(n6392), .ZN(n6002) );
  NAND4_X1 U5574 ( .A1(n5982), .A2(n5981), .A3(n5980), .A4(n5979), .ZN(n5983)
         );
  AOI22_X1 U5575 ( .A1(n4812), .A2(reg_file[520]), .B1(n4809), .B2(
        reg_file[552]), .ZN(n5979) );
  AOI22_X1 U5576 ( .A1(n3285), .A2(reg_file[616]), .B1(n4804), .B2(
        reg_file[584]), .ZN(n5980) );
  AOI22_X1 U5577 ( .A1(n3356), .A2(reg_file[712]), .B1(n4794), .B2(
        reg_file[680]), .ZN(n5981) );
  AOI22_X1 U5578 ( .A1(n4790), .A2(reg_file[648]), .B1(n4815), .B2(
        reg_file[744]), .ZN(n5982) );
  NAND2_X1 U5579 ( .A1(n5335), .A2(n3361), .ZN(n5336) );
  NAND4_X1 U5580 ( .A1(n5334), .A2(n5333), .A3(n5332), .A4(n5331), .ZN(n5335)
         );
  AOI22_X1 U5581 ( .A1(n3296), .A2(reg_file[776]), .B1(n3318), .B2(
        reg_file[808]), .ZN(n5331) );
  AOI22_X1 U5582 ( .A1(n4784), .A2(reg_file[872]), .B1(n4771), .B2(
        reg_file[840]), .ZN(n5332) );
  AOI22_X1 U5583 ( .A1(n3294), .A2(reg_file[936]), .B1(n4763), .B2(
        reg_file[904]), .ZN(n5333) );
  AOI22_X1 U5584 ( .A1(n4756), .A2(reg_file[968]), .B1(n4759), .B2(
        reg_file[1000]), .ZN(n5334) );
  NAND2_X1 U5585 ( .A1(n5330), .A2(n3390), .ZN(n5337) );
  NAND4_X1 U5586 ( .A1(n5329), .A2(n5328), .A3(n5327), .A4(n5326), .ZN(n5330)
         );
  AOI22_X1 U5587 ( .A1(n3296), .A2(reg_file[520]), .B1(n3318), .B2(
        reg_file[552]), .ZN(n5326) );
  AOI22_X1 U5588 ( .A1(n4784), .A2(reg_file[616]), .B1(n4771), .B2(
        reg_file[584]), .ZN(n5327) );
  AOI22_X1 U5589 ( .A1(n3294), .A2(reg_file[680]), .B1(n4763), .B2(
        reg_file[648]), .ZN(n5328) );
  AOI22_X1 U5590 ( .A1(n4757), .A2(reg_file[712]), .B1(n4759), .B2(
        reg_file[744]), .ZN(n5329) );
  NAND2_X1 U5591 ( .A1(n5325), .A2(n5805), .ZN(n5338) );
  NAND4_X1 U5592 ( .A1(n5324), .A2(n5323), .A3(n5322), .A4(n5321), .ZN(n5325)
         );
  AOI22_X1 U5593 ( .A1(n3296), .A2(reg_file[8]), .B1(n3318), .B2(reg_file[40]), 
        .ZN(n5321) );
  AOI22_X1 U5594 ( .A1(n4784), .A2(reg_file[104]), .B1(n4771), .B2(
        reg_file[72]), .ZN(n5322) );
  AOI22_X1 U5595 ( .A1(n3294), .A2(reg_file[168]), .B1(n4763), .B2(
        reg_file[136]), .ZN(n5323) );
  AOI22_X1 U5596 ( .A1(n4757), .A2(reg_file[200]), .B1(n4759), .B2(
        reg_file[232]), .ZN(n5324) );
  NAND2_X1 U5597 ( .A1(n5320), .A2(n3389), .ZN(n5339) );
  NAND4_X1 U5598 ( .A1(n5319), .A2(n5318), .A3(n5317), .A4(n5316), .ZN(n5320)
         );
  AOI22_X1 U5599 ( .A1(n3296), .A2(reg_file[264]), .B1(n3318), .B2(
        reg_file[296]), .ZN(n5316) );
  AOI22_X1 U5600 ( .A1(n4784), .A2(reg_file[360]), .B1(n4771), .B2(
        reg_file[328]), .ZN(n5317) );
  AOI22_X1 U5601 ( .A1(n3294), .A2(reg_file[424]), .B1(n4763), .B2(
        reg_file[392]), .ZN(n5318) );
  AOI22_X1 U5602 ( .A1(n5809), .A2(reg_file[456]), .B1(n4759), .B2(
        reg_file[488]), .ZN(n5319) );
  NAND2_X1 U5603 ( .A1(n5950), .A2(n3362), .ZN(n5951) );
  NAND4_X1 U5604 ( .A1(n5949), .A2(n5948), .A3(n5947), .A4(n5946), .ZN(n5950)
         );
  AOI22_X1 U5605 ( .A1(n4812), .A2(reg_file[774]), .B1(n4808), .B2(
        reg_file[806]), .ZN(n5946) );
  AOI22_X1 U5606 ( .A1(n3286), .A2(reg_file[870]), .B1(n4804), .B2(
        reg_file[838]), .ZN(n5947) );
  AOI22_X1 U5607 ( .A1(n4800), .A2(reg_file[966]), .B1(n4797), .B2(
        reg_file[934]), .ZN(n5948) );
  AOI22_X1 U5608 ( .A1(reg_file[902]), .A2(n3386), .B1(n4815), .B2(
        reg_file[998]), .ZN(n5949) );
  NAND2_X1 U5609 ( .A1(n5945), .A2(n6392), .ZN(n5952) );
  NAND4_X1 U5610 ( .A1(n5944), .A2(n5943), .A3(n5942), .A4(n5941), .ZN(n5945)
         );
  AOI22_X1 U5611 ( .A1(n4811), .A2(reg_file[518]), .B1(n4807), .B2(
        reg_file[550]), .ZN(n5941) );
  AOI22_X1 U5612 ( .A1(n3286), .A2(reg_file[614]), .B1(n4804), .B2(
        reg_file[582]), .ZN(n5942) );
  AOI22_X1 U5613 ( .A1(n4801), .A2(reg_file[710]), .B1(n4797), .B2(
        reg_file[678]), .ZN(n5943) );
  AOI22_X1 U5614 ( .A1(n3355), .A2(reg_file[646]), .B1(n4815), .B2(
        reg_file[742]), .ZN(n5944) );
  NAND2_X1 U5615 ( .A1(n5940), .A2(n6381), .ZN(n5953) );
  NAND4_X1 U5616 ( .A1(n5939), .A2(n5938), .A3(n5937), .A4(n5936), .ZN(n5940)
         );
  AOI22_X1 U5617 ( .A1(n4811), .A2(reg_file[262]), .B1(n4808), .B2(
        reg_file[294]), .ZN(n5936) );
  AOI22_X1 U5618 ( .A1(n3285), .A2(reg_file[358]), .B1(n4804), .B2(
        reg_file[326]), .ZN(n5937) );
  AOI22_X1 U5619 ( .A1(n4801), .A2(reg_file[454]), .B1(n4796), .B2(
        reg_file[422]), .ZN(n5938) );
  AOI22_X1 U5620 ( .A1(n3355), .A2(reg_file[390]), .B1(n4815), .B2(
        reg_file[486]), .ZN(n5939) );
  NAND2_X1 U5621 ( .A1(n5935), .A2(n6373), .ZN(n5954) );
  NAND4_X1 U5622 ( .A1(n5934), .A2(n5933), .A3(n5932), .A4(n5931), .ZN(n5935)
         );
  AOI22_X1 U5623 ( .A1(n4812), .A2(reg_file[6]), .B1(n4807), .B2(reg_file[38]), 
        .ZN(n5931) );
  AOI22_X1 U5624 ( .A1(n3286), .A2(reg_file[102]), .B1(n4804), .B2(
        reg_file[70]), .ZN(n5932) );
  AOI22_X1 U5625 ( .A1(n3356), .A2(reg_file[198]), .B1(n4795), .B2(
        reg_file[166]), .ZN(n5933) );
  AOI22_X1 U5626 ( .A1(n3355), .A2(reg_file[134]), .B1(n4815), .B2(
        reg_file[230]), .ZN(n5934) );
  NAND4_X1 U5627 ( .A1(n5291), .A2(n5290), .A3(n5289), .A4(n5288), .ZN(
        rs2_val_gpr_w[6]) );
  NAND2_X1 U5628 ( .A1(n5287), .A2(n3390), .ZN(n5288) );
  NAND4_X1 U5629 ( .A1(n5286), .A2(n5285), .A3(n5284), .A4(n5283), .ZN(n5287)
         );
  AOI22_X1 U5630 ( .A1(n3296), .A2(reg_file[518]), .B1(n3318), .B2(
        reg_file[550]), .ZN(n5283) );
  AOI22_X1 U5631 ( .A1(n4784), .A2(reg_file[614]), .B1(n4771), .B2(
        reg_file[582]), .ZN(n5284) );
  AOI22_X1 U5632 ( .A1(n3294), .A2(reg_file[678]), .B1(n4763), .B2(
        reg_file[646]), .ZN(n5285) );
  AOI22_X1 U5633 ( .A1(n4756), .A2(reg_file[710]), .B1(n4758), .B2(
        reg_file[742]), .ZN(n5286) );
  NAND2_X1 U5634 ( .A1(n5282), .A2(n5805), .ZN(n5289) );
  NAND4_X1 U5635 ( .A1(n5281), .A2(n5280), .A3(n5279), .A4(n5278), .ZN(n5282)
         );
  AOI22_X1 U5636 ( .A1(n3296), .A2(reg_file[6]), .B1(n3318), .B2(reg_file[38]), 
        .ZN(n5278) );
  AOI22_X1 U5637 ( .A1(n4784), .A2(reg_file[102]), .B1(n4771), .B2(
        reg_file[70]), .ZN(n5279) );
  AOI22_X1 U5638 ( .A1(n3294), .A2(reg_file[166]), .B1(n4763), .B2(
        reg_file[134]), .ZN(n5280) );
  AOI22_X1 U5639 ( .A1(n3519), .A2(reg_file[198]), .B1(n4758), .B2(
        reg_file[230]), .ZN(n5281) );
  NAND2_X1 U5640 ( .A1(n5277), .A2(n3361), .ZN(n5290) );
  NAND4_X1 U5641 ( .A1(n5276), .A2(n5275), .A3(n5274), .A4(n5273), .ZN(n5277)
         );
  AOI22_X1 U5642 ( .A1(n3296), .A2(reg_file[774]), .B1(n3318), .B2(
        reg_file[806]), .ZN(n5273) );
  AOI22_X1 U5643 ( .A1(n4784), .A2(reg_file[870]), .B1(n4771), .B2(
        reg_file[838]), .ZN(n5274) );
  AOI22_X1 U5644 ( .A1(n3294), .A2(reg_file[934]), .B1(n4763), .B2(
        reg_file[902]), .ZN(n5275) );
  AOI22_X1 U5645 ( .A1(n4757), .A2(reg_file[966]), .B1(n4758), .B2(
        reg_file[998]), .ZN(n5276) );
  NAND2_X1 U5646 ( .A1(n5272), .A2(n3389), .ZN(n5291) );
  NAND4_X1 U5647 ( .A1(n5271), .A2(n5270), .A3(n5269), .A4(n5268), .ZN(n5272)
         );
  AOI22_X1 U5648 ( .A1(n3296), .A2(reg_file[262]), .B1(n3318), .B2(
        reg_file[294]), .ZN(n5268) );
  AOI22_X1 U5649 ( .A1(n4784), .A2(reg_file[358]), .B1(n4771), .B2(
        reg_file[326]), .ZN(n5269) );
  AOI22_X1 U5650 ( .A1(n3294), .A2(reg_file[422]), .B1(n4763), .B2(
        reg_file[390]), .ZN(n5270) );
  AOI22_X1 U5651 ( .A1(n4756), .A2(reg_file[454]), .B1(n4758), .B2(
        reg_file[486]), .ZN(n5271) );
  NAND2_X1 U5652 ( .A1(n5974), .A2(n3362), .ZN(n5975) );
  NAND4_X1 U5653 ( .A1(n5973), .A2(n5972), .A3(n5971), .A4(n5970), .ZN(n5974)
         );
  AOI22_X1 U5654 ( .A1(n4811), .A2(reg_file[775]), .B1(n4808), .B2(
        reg_file[807]), .ZN(n5970) );
  AOI22_X1 U5655 ( .A1(n3285), .A2(reg_file[871]), .B1(n4804), .B2(
        reg_file[839]), .ZN(n5971) );
  AOI22_X1 U5656 ( .A1(n4799), .A2(reg_file[967]), .B1(n3360), .B2(
        reg_file[935]), .ZN(n5972) );
  AOI22_X1 U5657 ( .A1(n3355), .A2(reg_file[903]), .B1(n4815), .B2(
        reg_file[999]), .ZN(n5973) );
  NAND2_X1 U5658 ( .A1(n5969), .A2(n6392), .ZN(n5976) );
  NAND4_X1 U5659 ( .A1(n5968), .A2(n5967), .A3(n5966), .A4(n5965), .ZN(n5969)
         );
  AOI22_X1 U5660 ( .A1(n4812), .A2(reg_file[519]), .B1(n4809), .B2(
        reg_file[551]), .ZN(n5965) );
  AOI22_X1 U5661 ( .A1(n3285), .A2(reg_file[615]), .B1(n4804), .B2(
        reg_file[583]), .ZN(n5966) );
  AOI22_X1 U5662 ( .A1(n4801), .A2(reg_file[711]), .B1(n3360), .B2(
        reg_file[679]), .ZN(n5967) );
  AOI22_X1 U5663 ( .A1(n3355), .A2(reg_file[647]), .B1(n4815), .B2(
        reg_file[743]), .ZN(n5968) );
  NAND2_X1 U5664 ( .A1(n5964), .A2(n6381), .ZN(n5977) );
  NAND4_X1 U5665 ( .A1(n5963), .A2(n5962), .A3(n5961), .A4(n5960), .ZN(n5964)
         );
  AOI22_X1 U5666 ( .A1(n4811), .A2(reg_file[263]), .B1(n4807), .B2(
        reg_file[295]), .ZN(n5960) );
  AOI22_X1 U5667 ( .A1(n3285), .A2(reg_file[359]), .B1(n4804), .B2(
        reg_file[327]), .ZN(n5961) );
  AOI22_X1 U5668 ( .A1(n4798), .A2(reg_file[455]), .B1(n4795), .B2(
        reg_file[423]), .ZN(n5962) );
  AOI22_X1 U5669 ( .A1(reg_file[391]), .A2(n3355), .B1(n4815), .B2(
        reg_file[487]), .ZN(n5963) );
  NAND2_X1 U5670 ( .A1(n5959), .A2(n6373), .ZN(n5978) );
  NAND4_X1 U5671 ( .A1(n5958), .A2(n5957), .A3(n5956), .A4(n5955), .ZN(n5959)
         );
  AOI22_X1 U5672 ( .A1(n4812), .A2(reg_file[7]), .B1(n4809), .B2(reg_file[39]), 
        .ZN(n5955) );
  AOI22_X1 U5673 ( .A1(n3285), .A2(reg_file[103]), .B1(n4804), .B2(
        reg_file[71]), .ZN(n5956) );
  AOI22_X1 U5674 ( .A1(n4800), .A2(reg_file[199]), .B1(n4796), .B2(
        reg_file[167]), .ZN(n5957) );
  AOI22_X1 U5675 ( .A1(reg_file[135]), .A2(n3355), .B1(n4815), .B2(
        reg_file[231]), .ZN(n5958) );
  NAND2_X1 U5676 ( .A1(n5311), .A2(n3390), .ZN(n5312) );
  NAND4_X1 U5677 ( .A1(n5310), .A2(n5309), .A3(n5308), .A4(n5307), .ZN(n5311)
         );
  AOI22_X1 U5678 ( .A1(n3296), .A2(reg_file[519]), .B1(n3318), .B2(
        reg_file[551]), .ZN(n5307) );
  AOI22_X1 U5679 ( .A1(n4784), .A2(reg_file[615]), .B1(n4771), .B2(
        reg_file[583]), .ZN(n5308) );
  AOI22_X1 U5680 ( .A1(n3294), .A2(reg_file[679]), .B1(n4763), .B2(
        reg_file[647]), .ZN(n5309) );
  AOI22_X1 U5681 ( .A1(n4757), .A2(reg_file[711]), .B1(n4759), .B2(
        reg_file[743]), .ZN(n5310) );
  NAND2_X1 U5682 ( .A1(n5306), .A2(n5805), .ZN(n5313) );
  NAND4_X1 U5683 ( .A1(n5305), .A2(n5304), .A3(n5303), .A4(n5302), .ZN(n5306)
         );
  AOI22_X1 U5684 ( .A1(n3296), .A2(reg_file[7]), .B1(n3318), .B2(reg_file[39]), 
        .ZN(n5302) );
  AOI22_X1 U5685 ( .A1(n4784), .A2(reg_file[103]), .B1(n4771), .B2(
        reg_file[71]), .ZN(n5303) );
  AOI22_X1 U5686 ( .A1(n3294), .A2(reg_file[167]), .B1(n4763), .B2(
        reg_file[135]), .ZN(n5304) );
  AOI22_X1 U5687 ( .A1(n4757), .A2(reg_file[199]), .B1(n4759), .B2(
        reg_file[231]), .ZN(n5305) );
  NAND2_X1 U5688 ( .A1(n5301), .A2(n3361), .ZN(n5314) );
  NAND4_X1 U5689 ( .A1(n5300), .A2(n5299), .A3(n5298), .A4(n5297), .ZN(n5301)
         );
  AOI22_X1 U5690 ( .A1(n3296), .A2(reg_file[775]), .B1(n3318), .B2(
        reg_file[807]), .ZN(n5297) );
  AOI22_X1 U5691 ( .A1(n4784), .A2(reg_file[871]), .B1(n4771), .B2(
        reg_file[839]), .ZN(n5298) );
  AOI22_X1 U5692 ( .A1(n3294), .A2(reg_file[935]), .B1(n4763), .B2(
        reg_file[903]), .ZN(n5299) );
  AOI22_X1 U5693 ( .A1(n4755), .A2(reg_file[967]), .B1(n4759), .B2(
        reg_file[999]), .ZN(n5300) );
  NAND2_X1 U5694 ( .A1(n5296), .A2(n3389), .ZN(n5315) );
  NAND4_X1 U5695 ( .A1(n5295), .A2(n5294), .A3(n5293), .A4(n5292), .ZN(n5296)
         );
  AOI22_X1 U5696 ( .A1(n3296), .A2(reg_file[263]), .B1(n3318), .B2(
        reg_file[295]), .ZN(n5292) );
  AOI22_X1 U5697 ( .A1(n4784), .A2(reg_file[359]), .B1(n4771), .B2(
        reg_file[327]), .ZN(n5293) );
  AOI22_X1 U5698 ( .A1(n3294), .A2(reg_file[423]), .B1(n4763), .B2(
        reg_file[391]), .ZN(n5294) );
  AOI22_X1 U5699 ( .A1(n4757), .A2(reg_file[455]), .B1(n4759), .B2(
        reg_file[487]), .ZN(n5295) );
  NAND2_X1 U5700 ( .A1(n6022), .A2(n3362), .ZN(n6023) );
  NAND4_X1 U5701 ( .A1(n6021), .A2(n6020), .A3(n6019), .A4(n6018), .ZN(n6022)
         );
  AOI22_X1 U5702 ( .A1(n4812), .A2(reg_file[777]), .B1(n4808), .B2(
        reg_file[809]), .ZN(n6018) );
  AOI22_X1 U5703 ( .A1(n3286), .A2(reg_file[873]), .B1(n3295), .B2(
        reg_file[841]), .ZN(n6019) );
  AOI22_X1 U5704 ( .A1(n4799), .A2(reg_file[969]), .B1(n4792), .B2(
        reg_file[937]), .ZN(n6020) );
  AOI22_X1 U5705 ( .A1(n3355), .A2(reg_file[905]), .B1(n4815), .B2(
        reg_file[1001]), .ZN(n6021) );
  NAND2_X1 U5706 ( .A1(n6017), .A2(n6373), .ZN(n6024) );
  NAND4_X1 U5707 ( .A1(n6016), .A2(n6015), .A3(n6014), .A4(n6013), .ZN(n6017)
         );
  AOI22_X1 U5708 ( .A1(n4812), .A2(reg_file[9]), .B1(n4808), .B2(reg_file[41]), 
        .ZN(n6013) );
  AOI22_X1 U5709 ( .A1(n3285), .A2(reg_file[105]), .B1(n3295), .B2(
        reg_file[73]), .ZN(n6014) );
  AOI22_X1 U5710 ( .A1(n4799), .A2(reg_file[201]), .B1(n4792), .B2(
        reg_file[169]), .ZN(n6015) );
  AOI22_X1 U5711 ( .A1(n3355), .A2(reg_file[137]), .B1(n4815), .B2(
        reg_file[233]), .ZN(n6016) );
  NAND2_X1 U5712 ( .A1(n6012), .A2(n6381), .ZN(n6025) );
  NAND4_X1 U5713 ( .A1(n6011), .A2(n6010), .A3(n6009), .A4(n6008), .ZN(n6012)
         );
  AOI22_X1 U5714 ( .A1(n4812), .A2(reg_file[265]), .B1(n4808), .B2(
        reg_file[297]), .ZN(n6008) );
  AOI22_X1 U5715 ( .A1(n3286), .A2(reg_file[361]), .B1(n3295), .B2(
        reg_file[329]), .ZN(n6009) );
  AOI22_X1 U5716 ( .A1(n4799), .A2(reg_file[457]), .B1(n4792), .B2(
        reg_file[425]), .ZN(n6010) );
  AOI22_X1 U5717 ( .A1(reg_file[393]), .A2(n3386), .B1(n4815), .B2(
        reg_file[489]), .ZN(n6011) );
  NAND2_X1 U5718 ( .A1(n6007), .A2(n6392), .ZN(n6026) );
  NAND4_X1 U5719 ( .A1(n6006), .A2(n6005), .A3(n6004), .A4(n6003), .ZN(n6007)
         );
  AOI22_X1 U5720 ( .A1(n4812), .A2(reg_file[521]), .B1(n4808), .B2(
        reg_file[553]), .ZN(n6003) );
  AOI22_X1 U5721 ( .A1(n3286), .A2(reg_file[617]), .B1(n3295), .B2(
        reg_file[585]), .ZN(n6004) );
  AOI22_X1 U5722 ( .A1(n4799), .A2(reg_file[713]), .B1(n4792), .B2(
        reg_file[681]), .ZN(n6005) );
  AOI22_X1 U5723 ( .A1(n3386), .A2(reg_file[649]), .B1(n4815), .B2(
        reg_file[745]), .ZN(n6006) );
  NAND2_X1 U5724 ( .A1(n5359), .A2(n3361), .ZN(n5360) );
  NAND4_X1 U5725 ( .A1(n5358), .A2(n5357), .A3(n5356), .A4(n5355), .ZN(n5359)
         );
  AOI22_X1 U5726 ( .A1(n4789), .A2(reg_file[777]), .B1(n4786), .B2(
        reg_file[809]), .ZN(n5355) );
  AOI22_X1 U5727 ( .A1(n4783), .A2(reg_file[873]), .B1(n4772), .B2(
        reg_file[841]), .ZN(n5356) );
  AOI22_X1 U5728 ( .A1(n3294), .A2(reg_file[937]), .B1(n4767), .B2(
        reg_file[905]), .ZN(n5357) );
  AOI22_X1 U5729 ( .A1(n3519), .A2(reg_file[969]), .B1(n4759), .B2(
        reg_file[1001]), .ZN(n5358) );
  NAND2_X1 U5730 ( .A1(n5354), .A2(n5805), .ZN(n5361) );
  NAND4_X1 U5731 ( .A1(n5353), .A2(n5352), .A3(n5351), .A4(n5350), .ZN(n5354)
         );
  AOI22_X1 U5732 ( .A1(n4789), .A2(reg_file[9]), .B1(n4787), .B2(reg_file[41]), 
        .ZN(n5350) );
  AOI22_X1 U5733 ( .A1(n4783), .A2(reg_file[105]), .B1(n4772), .B2(
        reg_file[73]), .ZN(n5351) );
  AOI22_X1 U5734 ( .A1(n3294), .A2(reg_file[169]), .B1(n4768), .B2(
        reg_file[137]), .ZN(n5352) );
  AOI22_X1 U5735 ( .A1(n4756), .A2(reg_file[201]), .B1(n4759), .B2(
        reg_file[233]), .ZN(n5353) );
  NAND2_X1 U5736 ( .A1(n5349), .A2(n3390), .ZN(n5362) );
  NAND4_X1 U5737 ( .A1(n5348), .A2(n5347), .A3(n5346), .A4(n5345), .ZN(n5349)
         );
  AOI22_X1 U5738 ( .A1(n4789), .A2(reg_file[521]), .B1(n4786), .B2(
        reg_file[553]), .ZN(n5345) );
  AOI22_X1 U5739 ( .A1(n4783), .A2(reg_file[617]), .B1(n4772), .B2(
        reg_file[585]), .ZN(n5346) );
  AOI22_X1 U5740 ( .A1(n3294), .A2(reg_file[681]), .B1(n4768), .B2(
        reg_file[649]), .ZN(n5347) );
  AOI22_X1 U5741 ( .A1(n4757), .A2(reg_file[713]), .B1(n4759), .B2(
        reg_file[745]), .ZN(n5348) );
  NAND2_X1 U5742 ( .A1(n5344), .A2(n3389), .ZN(n5363) );
  NAND4_X1 U5743 ( .A1(n5343), .A2(n5342), .A3(n5341), .A4(n5340), .ZN(n5344)
         );
  AOI22_X1 U5744 ( .A1(n3296), .A2(reg_file[265]), .B1(n4787), .B2(
        reg_file[297]), .ZN(n5340) );
  AOI22_X1 U5745 ( .A1(n4784), .A2(reg_file[361]), .B1(n4772), .B2(
        reg_file[329]), .ZN(n5341) );
  AOI22_X1 U5746 ( .A1(n3294), .A2(reg_file[425]), .B1(n3769), .B2(
        reg_file[393]), .ZN(n5342) );
  AOI22_X1 U5747 ( .A1(n4755), .A2(reg_file[457]), .B1(n4759), .B2(
        reg_file[489]), .ZN(n5343) );
  AOI22_X1 U5748 ( .A1(n4811), .A2(reg_file[517]), .B1(n4807), .B2(
        reg_file[549]), .ZN(n5927) );
  AOI22_X1 U5749 ( .A1(n3286), .A2(reg_file[613]), .B1(n4803), .B2(
        reg_file[581]), .ZN(n5928) );
  AOI22_X1 U5750 ( .A1(n4800), .A2(reg_file[709]), .B1(n4791), .B2(
        reg_file[677]), .ZN(n5929) );
  AOI22_X1 U5751 ( .A1(n3355), .A2(reg_file[645]), .B1(n3293), .B2(
        reg_file[741]), .ZN(n5930) );
  NAND4_X1 U5752 ( .A1(n5925), .A2(n5924), .A3(n5923), .A4(n5922), .ZN(n5926)
         );
  AOI22_X1 U5753 ( .A1(n4811), .A2(reg_file[5]), .B1(n4807), .B2(reg_file[37]), 
        .ZN(n5922) );
  AOI22_X1 U5754 ( .A1(n3285), .A2(reg_file[101]), .B1(n4803), .B2(
        reg_file[69]), .ZN(n5923) );
  AOI22_X1 U5755 ( .A1(n4801), .A2(reg_file[197]), .B1(n4791), .B2(
        reg_file[165]), .ZN(n5924) );
  AOI22_X1 U5756 ( .A1(n3355), .A2(reg_file[133]), .B1(n3293), .B2(
        reg_file[229]), .ZN(n5925) );
  AOI22_X1 U5757 ( .A1(n4811), .A2(reg_file[773]), .B1(n4807), .B2(
        reg_file[805]), .ZN(n5918) );
  AOI22_X1 U5758 ( .A1(n3285), .A2(reg_file[869]), .B1(n4803), .B2(
        reg_file[837]), .ZN(n5919) );
  AOI22_X1 U5759 ( .A1(n4801), .A2(reg_file[965]), .B1(n4791), .B2(
        reg_file[933]), .ZN(n5920) );
  AOI22_X1 U5760 ( .A1(n4790), .A2(reg_file[901]), .B1(n3354), .B2(
        reg_file[997]), .ZN(n5921) );
  AOI22_X1 U5761 ( .A1(n4811), .A2(reg_file[261]), .B1(n4807), .B2(
        reg_file[293]), .ZN(n5914) );
  AOI22_X1 U5762 ( .A1(n3285), .A2(reg_file[357]), .B1(n4803), .B2(
        reg_file[325]), .ZN(n5915) );
  AOI22_X1 U5763 ( .A1(n4801), .A2(reg_file[453]), .B1(n4791), .B2(
        reg_file[421]), .ZN(n5916) );
  AOI22_X1 U5764 ( .A1(n3355), .A2(reg_file[389]), .B1(n3293), .B2(
        reg_file[485]), .ZN(n5917) );
  AOI22_X1 U5765 ( .A1(n4788), .A2(reg_file[517]), .B1(n3318), .B2(
        reg_file[549]), .ZN(n5264) );
  AOI22_X1 U5766 ( .A1(n4785), .A2(reg_file[613]), .B1(n4770), .B2(
        reg_file[581]), .ZN(n5265) );
  AOI22_X1 U5767 ( .A1(n3357), .A2(reg_file[677]), .B1(n4762), .B2(
        reg_file[645]), .ZN(n5266) );
  AOI22_X1 U5768 ( .A1(n4757), .A2(reg_file[709]), .B1(n4760), .B2(
        reg_file[741]), .ZN(n5267) );
  AOI22_X1 U5769 ( .A1(n4788), .A2(reg_file[261]), .B1(n3318), .B2(
        reg_file[293]), .ZN(n5260) );
  AOI22_X1 U5770 ( .A1(n4785), .A2(reg_file[357]), .B1(n4770), .B2(
        reg_file[325]), .ZN(n5261) );
  AOI22_X1 U5771 ( .A1(n3357), .A2(reg_file[421]), .B1(n4762), .B2(
        reg_file[389]), .ZN(n5262) );
  AOI22_X1 U5772 ( .A1(n4756), .A2(reg_file[453]), .B1(n4760), .B2(
        reg_file[485]), .ZN(n5263) );
  AOI22_X1 U5773 ( .A1(n4788), .A2(reg_file[773]), .B1(n3318), .B2(
        reg_file[805]), .ZN(n5256) );
  AOI22_X1 U5774 ( .A1(n4785), .A2(reg_file[869]), .B1(n4770), .B2(
        reg_file[837]), .ZN(n5257) );
  AOI22_X1 U5775 ( .A1(n3357), .A2(reg_file[933]), .B1(n4762), .B2(
        reg_file[901]), .ZN(n5258) );
  AOI22_X1 U5776 ( .A1(n4757), .A2(reg_file[965]), .B1(n4760), .B2(
        reg_file[997]), .ZN(n5259) );
  AOI22_X1 U5777 ( .A1(n4788), .A2(reg_file[5]), .B1(n3318), .B2(reg_file[37]), 
        .ZN(n5253) );
  AOI22_X1 U5778 ( .A1(n4785), .A2(reg_file[101]), .B1(n4770), .B2(
        reg_file[69]), .ZN(n5254) );
  AOI22_X1 U5779 ( .A1(n3357), .A2(reg_file[165]), .B1(n4762), .B2(
        reg_file[133]), .ZN(n5255) );
  NAND2_X1 U5780 ( .A1(n5053), .A2(n3390), .ZN(n5054) );
  NAND4_X1 U5781 ( .A1(n5052), .A2(n5051), .A3(n5050), .A4(n5049), .ZN(n5053)
         );
  AOI22_X1 U5782 ( .A1(n5809), .A2(reg_file[705]), .B1(n5810), .B2(
        reg_file[737]), .ZN(n5052) );
  NAND2_X1 U5783 ( .A1(n5048), .A2(n3389), .ZN(n5055) );
  NAND4_X1 U5784 ( .A1(n5047), .A2(n5046), .A3(n5045), .A4(n5044), .ZN(n5048)
         );
  AOI22_X1 U5785 ( .A1(n4756), .A2(reg_file[449]), .B1(n5810), .B2(
        reg_file[481]), .ZN(n5047) );
  NAND2_X1 U5786 ( .A1(n5043), .A2(n3361), .ZN(n5056) );
  NAND4_X1 U5787 ( .A1(n5042), .A2(n5041), .A3(n5040), .A4(n5039), .ZN(n5043)
         );
  AOI22_X1 U5788 ( .A1(n4756), .A2(reg_file[961]), .B1(n5810), .B2(
        reg_file[993]), .ZN(n5042) );
  NAND2_X1 U5789 ( .A1(n5038), .A2(n5805), .ZN(n5057) );
  NAND4_X1 U5790 ( .A1(n5037), .A2(n5036), .A3(n5035), .A4(n5034), .ZN(n5038)
         );
  AOI22_X1 U5791 ( .A1(n4756), .A2(reg_file[193]), .B1(n5810), .B2(
        reg_file[225]), .ZN(n5037) );
  NAND2_X1 U5792 ( .A1(n4996), .A2(n3361), .ZN(n4997) );
  NAND4_X1 U5793 ( .A1(n4995), .A2(n4994), .A3(n4993), .A4(n4992), .ZN(n4996)
         );
  AOI22_X1 U5794 ( .A1(n3519), .A2(reg_file[960]), .B1(n5810), .B2(
        reg_file[992]), .ZN(n4995) );
  NAND2_X1 U5795 ( .A1(n4991), .A2(n5805), .ZN(n4998) );
  NAND4_X1 U5796 ( .A1(n4990), .A2(n4989), .A3(n4988), .A4(n4987), .ZN(n4991)
         );
  AOI22_X1 U5797 ( .A1(n3519), .A2(reg_file[192]), .B1(n5810), .B2(
        reg_file[224]), .ZN(n4990) );
  NAND2_X1 U5798 ( .A1(n4986), .A2(n3390), .ZN(n4999) );
  NAND4_X1 U5799 ( .A1(n4985), .A2(n4984), .A3(n4983), .A4(n4982), .ZN(n4986)
         );
  AOI22_X1 U5800 ( .A1(n3519), .A2(reg_file[704]), .B1(n5810), .B2(
        reg_file[736]), .ZN(n4985) );
  NAND2_X1 U5801 ( .A1(n4981), .A2(n3389), .ZN(n5000) );
  NAND4_X1 U5802 ( .A1(n4980), .A2(n4979), .A3(n4978), .A4(n4977), .ZN(n4981)
         );
  AOI22_X1 U5803 ( .A1(n4755), .A2(reg_file[448]), .B1(n5810), .B2(
        reg_file[480]), .ZN(n4980) );
  NAND2_X1 U5804 ( .A1(n5861), .A2(n6392), .ZN(n5862) );
  NAND4_X1 U5805 ( .A1(n5859), .A2(n5860), .A3(n5858), .A4(n5857), .ZN(n5861)
         );
  NAND2_X1 U5806 ( .A1(n5856), .A2(n6373), .ZN(n5863) );
  NAND4_X1 U5807 ( .A1(n5855), .A2(n5854), .A3(n5853), .A4(n5852), .ZN(n5856)
         );
  NAND2_X1 U5808 ( .A1(n5851), .A2(n3362), .ZN(n5864) );
  NAND4_X1 U5809 ( .A1(n5850), .A2(n5849), .A3(n5848), .A4(n5847), .ZN(n5851)
         );
  NAND2_X1 U5810 ( .A1(n5846), .A2(n6381), .ZN(n5865) );
  NAND4_X1 U5811 ( .A1(n5845), .A2(n5844), .A3(n5843), .A4(n5842), .ZN(n5846)
         );
  NAND2_X1 U5812 ( .A1(n5110), .A2(n3361), .ZN(n5111) );
  NAND4_X1 U5813 ( .A1(n5109), .A2(n5108), .A3(n5107), .A4(n5106), .ZN(n5110)
         );
  AOI22_X1 U5814 ( .A1(n3519), .A2(reg_file[962]), .B1(n4760), .B2(
        reg_file[994]), .ZN(n5109) );
  NAND2_X1 U5815 ( .A1(n5105), .A2(n3389), .ZN(n5112) );
  NAND4_X1 U5816 ( .A1(n5104), .A2(n5103), .A3(n5102), .A4(n5101), .ZN(n5105)
         );
  AOI22_X1 U5817 ( .A1(n4755), .A2(reg_file[450]), .B1(n5810), .B2(
        reg_file[482]), .ZN(n5104) );
  NAND2_X1 U5818 ( .A1(n5100), .A2(n3390), .ZN(n5113) );
  NAND4_X1 U5819 ( .A1(n5099), .A2(n5098), .A3(n5097), .A4(n5096), .ZN(n5100)
         );
  AOI22_X1 U5820 ( .A1(n3519), .A2(reg_file[706]), .B1(n5810), .B2(
        reg_file[738]), .ZN(n5099) );
  NAND2_X1 U5821 ( .A1(n5095), .A2(n5805), .ZN(n5114) );
  NAND4_X1 U5822 ( .A1(n5094), .A2(n5093), .A3(n5092), .A4(n5091), .ZN(n5095)
         );
  AOI22_X1 U5823 ( .A1(n3519), .A2(reg_file[194]), .B1(n5810), .B2(
        reg_file[226]), .ZN(n5094) );
  NAND2_X1 U5824 ( .A1(n5885), .A2(n3362), .ZN(n5886) );
  NAND4_X1 U5825 ( .A1(n5884), .A2(n5883), .A3(n5882), .A4(n5881), .ZN(n5885)
         );
  AOI22_X1 U5826 ( .A1(n4811), .A2(reg_file[771]), .B1(n4807), .B2(
        reg_file[803]), .ZN(n5881) );
  AOI22_X1 U5827 ( .A1(n3285), .A2(reg_file[867]), .B1(n4803), .B2(
        reg_file[835]), .ZN(n5882) );
  AOI22_X1 U5828 ( .A1(n4800), .A2(reg_file[963]), .B1(n4791), .B2(
        reg_file[931]), .ZN(n5883) );
  AOI22_X1 U5829 ( .A1(n4790), .A2(reg_file[899]), .B1(n3354), .B2(
        reg_file[995]), .ZN(n5884) );
  NAND2_X1 U5830 ( .A1(n5880), .A2(n6392), .ZN(n5887) );
  NAND4_X1 U5831 ( .A1(n5879), .A2(n5878), .A3(n5877), .A4(n5876), .ZN(n5880)
         );
  AOI22_X1 U5832 ( .A1(n4811), .A2(reg_file[515]), .B1(n4807), .B2(
        reg_file[547]), .ZN(n5876) );
  AOI22_X1 U5833 ( .A1(n3285), .A2(reg_file[611]), .B1(n4803), .B2(
        reg_file[579]), .ZN(n5877) );
  AOI22_X1 U5834 ( .A1(n4800), .A2(reg_file[707]), .B1(n4791), .B2(
        reg_file[675]), .ZN(n5878) );
  AOI22_X1 U5835 ( .A1(n3355), .A2(reg_file[643]), .B1(n3354), .B2(
        reg_file[739]), .ZN(n5879) );
  NAND2_X1 U5836 ( .A1(n5875), .A2(n6381), .ZN(n5888) );
  NAND4_X1 U5837 ( .A1(n5874), .A2(n5873), .A3(n5872), .A4(n5871), .ZN(n5875)
         );
  AOI22_X1 U5838 ( .A1(n4811), .A2(reg_file[259]), .B1(n4807), .B2(
        reg_file[291]), .ZN(n5871) );
  AOI22_X1 U5839 ( .A1(n3285), .A2(reg_file[355]), .B1(n4803), .B2(
        reg_file[323]), .ZN(n5872) );
  AOI22_X1 U5840 ( .A1(n4801), .A2(reg_file[451]), .B1(n4791), .B2(
        reg_file[419]), .ZN(n5873) );
  AOI22_X1 U5841 ( .A1(reg_file[387]), .A2(n3355), .B1(n3354), .B2(
        reg_file[483]), .ZN(n5874) );
  NAND2_X1 U5842 ( .A1(n5870), .A2(n6373), .ZN(n5889) );
  NAND4_X1 U5843 ( .A1(n5869), .A2(n5868), .A3(n5867), .A4(n5866), .ZN(n5870)
         );
  AOI22_X1 U5844 ( .A1(n4811), .A2(reg_file[3]), .B1(n4807), .B2(reg_file[35]), 
        .ZN(n5866) );
  AOI22_X1 U5845 ( .A1(n3286), .A2(reg_file[99]), .B1(n4803), .B2(reg_file[67]), .ZN(n5867) );
  AOI22_X1 U5846 ( .A1(n4800), .A2(reg_file[195]), .B1(n4791), .B2(
        reg_file[163]), .ZN(n5868) );
  AOI22_X1 U5847 ( .A1(n3355), .A2(reg_file[131]), .B1(n3354), .B2(
        reg_file[227]), .ZN(n5869) );
  NAND2_X1 U5848 ( .A1(n5166), .A2(n3361), .ZN(n5167) );
  NAND4_X1 U5849 ( .A1(n5165), .A2(n5164), .A3(n5163), .A4(n5162), .ZN(n5166)
         );
  AOI22_X1 U5850 ( .A1(n3296), .A2(reg_file[771]), .B1(n3318), .B2(
        reg_file[803]), .ZN(n5162) );
  AOI22_X1 U5851 ( .A1(n4785), .A2(reg_file[867]), .B1(n4770), .B2(
        reg_file[835]), .ZN(n5163) );
  AOI22_X1 U5852 ( .A1(n3357), .A2(reg_file[931]), .B1(n4762), .B2(
        reg_file[899]), .ZN(n5164) );
  AOI22_X1 U5853 ( .A1(n4756), .A2(reg_file[963]), .B1(n4760), .B2(
        reg_file[995]), .ZN(n5165) );
  NAND2_X1 U5854 ( .A1(n5161), .A2(n3389), .ZN(n5168) );
  NAND4_X1 U5855 ( .A1(n5160), .A2(n5159), .A3(n5158), .A4(n5157), .ZN(n5161)
         );
  AOI22_X1 U5856 ( .A1(n4789), .A2(reg_file[259]), .B1(n3318), .B2(
        reg_file[291]), .ZN(n5157) );
  AOI22_X1 U5857 ( .A1(n4785), .A2(reg_file[355]), .B1(n4770), .B2(
        reg_file[323]), .ZN(n5158) );
  AOI22_X1 U5858 ( .A1(n3357), .A2(reg_file[419]), .B1(n4762), .B2(
        reg_file[387]), .ZN(n5159) );
  AOI22_X1 U5859 ( .A1(n4756), .A2(reg_file[451]), .B1(n4760), .B2(
        reg_file[483]), .ZN(n5160) );
  NAND2_X1 U5860 ( .A1(n5156), .A2(n3390), .ZN(n5169) );
  NAND4_X1 U5861 ( .A1(n5155), .A2(n5154), .A3(n5153), .A4(n5152), .ZN(n5156)
         );
  AOI22_X1 U5862 ( .A1(n5813), .A2(reg_file[515]), .B1(n3318), .B2(
        reg_file[547]), .ZN(n5152) );
  AOI22_X1 U5863 ( .A1(n4785), .A2(reg_file[611]), .B1(n4770), .B2(
        reg_file[579]), .ZN(n5153) );
  AOI22_X1 U5864 ( .A1(n3357), .A2(reg_file[675]), .B1(n4762), .B2(
        reg_file[643]), .ZN(n5154) );
  AOI22_X1 U5865 ( .A1(n3519), .A2(reg_file[707]), .B1(n4760), .B2(
        reg_file[739]), .ZN(n5155) );
  NAND2_X1 U5866 ( .A1(n5151), .A2(n5805), .ZN(n5170) );
  NAND4_X1 U5867 ( .A1(n5150), .A2(n5149), .A3(n5148), .A4(n5147), .ZN(n5151)
         );
  AOI22_X1 U5868 ( .A1(n4788), .A2(reg_file[3]), .B1(n3318), .B2(reg_file[35]), 
        .ZN(n5147) );
  AOI22_X1 U5869 ( .A1(n4785), .A2(reg_file[99]), .B1(n4770), .B2(reg_file[67]), .ZN(n5148) );
  AOI22_X1 U5870 ( .A1(n3357), .A2(reg_file[163]), .B1(n4762), .B2(
        reg_file[131]), .ZN(n5149) );
  AOI22_X1 U5871 ( .A1(n4755), .A2(reg_file[195]), .B1(n4760), .B2(
        reg_file[227]), .ZN(n5150) );
  NAND2_X1 U5872 ( .A1(n5909), .A2(n3362), .ZN(n5910) );
  NAND4_X1 U5873 ( .A1(n5908), .A2(n5907), .A3(n5906), .A4(n5905), .ZN(n5909)
         );
  AOI22_X1 U5874 ( .A1(n4811), .A2(reg_file[772]), .B1(n4807), .B2(
        reg_file[804]), .ZN(n5905) );
  AOI22_X1 U5875 ( .A1(n3286), .A2(reg_file[868]), .B1(n4803), .B2(
        reg_file[836]), .ZN(n5906) );
  AOI22_X1 U5876 ( .A1(n4800), .A2(reg_file[964]), .B1(n4791), .B2(
        reg_file[932]), .ZN(n5907) );
  AOI22_X1 U5877 ( .A1(n3355), .A2(reg_file[900]), .B1(n3293), .B2(
        reg_file[996]), .ZN(n5908) );
  NAND2_X1 U5878 ( .A1(n5904), .A2(n6392), .ZN(n5911) );
  NAND4_X1 U5879 ( .A1(n5903), .A2(n5902), .A3(n5901), .A4(n5900), .ZN(n5904)
         );
  AOI22_X1 U5880 ( .A1(n4811), .A2(reg_file[516]), .B1(n4807), .B2(
        reg_file[548]), .ZN(n5900) );
  AOI22_X1 U5881 ( .A1(n3285), .A2(reg_file[612]), .B1(n4803), .B2(
        reg_file[580]), .ZN(n5901) );
  AOI22_X1 U5882 ( .A1(n4800), .A2(reg_file[708]), .B1(n4791), .B2(
        reg_file[676]), .ZN(n5902) );
  AOI22_X1 U5883 ( .A1(reg_file[644]), .A2(n3355), .B1(n3354), .B2(
        reg_file[740]), .ZN(n5903) );
  NAND2_X1 U5884 ( .A1(n5899), .A2(n6381), .ZN(n5912) );
  NAND4_X1 U5885 ( .A1(n5898), .A2(n5897), .A3(n5896), .A4(n5895), .ZN(n5899)
         );
  AOI22_X1 U5886 ( .A1(n4811), .A2(reg_file[260]), .B1(n4807), .B2(
        reg_file[292]), .ZN(n5895) );
  AOI22_X1 U5887 ( .A1(n3285), .A2(reg_file[356]), .B1(n4803), .B2(
        reg_file[324]), .ZN(n5896) );
  AOI22_X1 U5888 ( .A1(n4801), .A2(reg_file[452]), .B1(n4791), .B2(
        reg_file[420]), .ZN(n5897) );
  AOI22_X1 U5889 ( .A1(n4790), .A2(reg_file[388]), .B1(n3293), .B2(
        reg_file[484]), .ZN(n5898) );
  NAND2_X1 U5890 ( .A1(n5894), .A2(n6373), .ZN(n5913) );
  NAND4_X1 U5891 ( .A1(n5893), .A2(n5892), .A3(n5891), .A4(n5890), .ZN(n5894)
         );
  AOI22_X1 U5892 ( .A1(n4811), .A2(reg_file[4]), .B1(n4807), .B2(reg_file[36]), 
        .ZN(n5890) );
  AOI22_X1 U5893 ( .A1(n3286), .A2(reg_file[100]), .B1(n4803), .B2(
        reg_file[68]), .ZN(n5891) );
  AOI22_X1 U5894 ( .A1(n4800), .A2(reg_file[196]), .B1(n4791), .B2(
        reg_file[164]), .ZN(n5892) );
  AOI22_X1 U5895 ( .A1(reg_file[132]), .A2(n4790), .B1(n3293), .B2(
        reg_file[228]), .ZN(n5893) );
  NAND4_X1 U5896 ( .A1(n5219), .A2(n5218), .A3(n5217), .A4(n5216), .ZN(n5220)
         );
  AOI22_X1 U5897 ( .A1(n4788), .A2(reg_file[516]), .B1(n3318), .B2(
        reg_file[548]), .ZN(n5216) );
  AOI22_X1 U5898 ( .A1(n4785), .A2(reg_file[612]), .B1(n4770), .B2(
        reg_file[580]), .ZN(n5217) );
  AOI22_X1 U5899 ( .A1(n3357), .A2(reg_file[676]), .B1(n4762), .B2(
        reg_file[644]), .ZN(n5218) );
  AOI22_X1 U5900 ( .A1(n4756), .A2(reg_file[708]), .B1(n4760), .B2(
        reg_file[740]), .ZN(n5219) );
  AOI22_X1 U5901 ( .A1(n5813), .A2(reg_file[4]), .B1(n3318), .B2(reg_file[36]), 
        .ZN(n5212) );
  AOI22_X1 U5902 ( .A1(n4785), .A2(reg_file[100]), .B1(n4770), .B2(
        reg_file[68]), .ZN(n5213) );
  AOI22_X1 U5903 ( .A1(n3357), .A2(reg_file[164]), .B1(n4762), .B2(
        reg_file[132]), .ZN(n5214) );
  AOI22_X1 U5904 ( .A1(n4757), .A2(reg_file[196]), .B1(n4760), .B2(
        reg_file[228]), .ZN(n5215) );
  AOI22_X1 U5905 ( .A1(n5813), .A2(reg_file[772]), .B1(n3318), .B2(
        reg_file[804]), .ZN(n5208) );
  AOI22_X1 U5906 ( .A1(n4785), .A2(reg_file[868]), .B1(n4770), .B2(
        reg_file[836]), .ZN(n5209) );
  AOI22_X1 U5907 ( .A1(n3357), .A2(reg_file[932]), .B1(n4762), .B2(
        reg_file[900]), .ZN(n5210) );
  AOI22_X1 U5908 ( .A1(n4757), .A2(reg_file[964]), .B1(n4760), .B2(
        reg_file[996]), .ZN(n5211) );
  NAND4_X1 U5909 ( .A1(n5206), .A2(n5205), .A3(n5204), .A4(n5203), .ZN(n5207)
         );
  AOI22_X1 U5910 ( .A1(n4788), .A2(reg_file[260]), .B1(n3318), .B2(
        reg_file[292]), .ZN(n5203) );
  AOI22_X1 U5911 ( .A1(n4785), .A2(reg_file[356]), .B1(n4770), .B2(
        reg_file[324]), .ZN(n5204) );
  AOI22_X1 U5912 ( .A1(n3357), .A2(reg_file[420]), .B1(n4762), .B2(
        reg_file[388]), .ZN(n5205) );
  AOI22_X1 U5913 ( .A1(n3519), .A2(reg_file[452]), .B1(n4760), .B2(
        reg_file[484]), .ZN(n5206) );
  NAND4_X1 U5914 ( .A1(n5635), .A2(n5634), .A3(n5633), .A4(n5632), .ZN(
        rs2_val_gpr_w[22]) );
  NAND2_X1 U5915 ( .A1(n5631), .A2(n3361), .ZN(n5632) );
  NAND4_X1 U5916 ( .A1(n5630), .A2(n5629), .A3(n5628), .A4(n5627), .ZN(n5631)
         );
  AOI22_X1 U5917 ( .A1(n4788), .A2(reg_file[790]), .B1(n4786), .B2(
        reg_file[822]), .ZN(n5627) );
  AOI22_X1 U5918 ( .A1(n4780), .A2(reg_file[886]), .B1(n4776), .B2(
        reg_file[854]), .ZN(n5628) );
  AOI22_X1 U5919 ( .A1(n3294), .A2(reg_file[950]), .B1(n3769), .B2(
        reg_file[918]), .ZN(n5629) );
  AOI22_X1 U5920 ( .A1(n4757), .A2(reg_file[982]), .B1(n4759), .B2(
        reg_file[1014]), .ZN(n5630) );
  NAND2_X1 U5921 ( .A1(n5626), .A2(n4754), .ZN(n5633) );
  NAND4_X1 U5922 ( .A1(n5625), .A2(n5624), .A3(n5623), .A4(n5622), .ZN(n5626)
         );
  AOI22_X1 U5923 ( .A1(n4788), .A2(reg_file[22]), .B1(n4787), .B2(reg_file[54]), .ZN(n5622) );
  AOI22_X1 U5924 ( .A1(n4780), .A2(reg_file[118]), .B1(n4776), .B2(
        reg_file[86]), .ZN(n5623) );
  AOI22_X1 U5925 ( .A1(n3294), .A2(reg_file[182]), .B1(n3769), .B2(
        reg_file[150]), .ZN(n5624) );
  AOI22_X1 U5926 ( .A1(n4756), .A2(reg_file[214]), .B1(n4758), .B2(
        reg_file[246]), .ZN(n5625) );
  NAND2_X1 U5927 ( .A1(n5621), .A2(n3390), .ZN(n5634) );
  NAND4_X1 U5928 ( .A1(n5620), .A2(n5619), .A3(n5618), .A4(n5617), .ZN(n5621)
         );
  AOI22_X1 U5929 ( .A1(n4788), .A2(reg_file[534]), .B1(n4787), .B2(
        reg_file[566]), .ZN(n5617) );
  AOI22_X1 U5930 ( .A1(n4780), .A2(reg_file[630]), .B1(n4776), .B2(
        reg_file[598]), .ZN(n5618) );
  AOI22_X1 U5931 ( .A1(n3294), .A2(reg_file[694]), .B1(n3769), .B2(
        reg_file[662]), .ZN(n5619) );
  AOI22_X1 U5932 ( .A1(n4757), .A2(reg_file[726]), .B1(n4758), .B2(
        reg_file[758]), .ZN(n5620) );
  NAND2_X1 U5933 ( .A1(n5616), .A2(n3389), .ZN(n5635) );
  NAND4_X1 U5934 ( .A1(n5615), .A2(n5614), .A3(n5613), .A4(n5612), .ZN(n5616)
         );
  AOI22_X1 U5935 ( .A1(n4788), .A2(reg_file[278]), .B1(n4786), .B2(
        reg_file[310]), .ZN(n5612) );
  AOI22_X1 U5936 ( .A1(n4781), .A2(reg_file[374]), .B1(n4776), .B2(
        reg_file[342]), .ZN(n5613) );
  BUF_X1 U5937 ( .A(n5811), .Z(n4781) );
  AOI22_X1 U5938 ( .A1(n3294), .A2(reg_file[438]), .B1(n3769), .B2(
        reg_file[406]), .ZN(n5614) );
  AOI22_X1 U5939 ( .A1(n4757), .A2(reg_file[470]), .B1(n4758), .B2(
        reg_file[502]), .ZN(n5615) );
  NAND4_X1 U5940 ( .A1(n6297), .A2(n6296), .A3(n6295), .A4(n6294), .ZN(
        rs1_val_gpr_w[23]) );
  NAND2_X1 U5941 ( .A1(n6293), .A2(n3387), .ZN(n6294) );
  NAND4_X1 U5942 ( .A1(n6292), .A2(n6291), .A3(n6290), .A4(n6289), .ZN(n6293)
         );
  AOI22_X1 U5943 ( .A1(n3358), .A2(reg_file[279]), .B1(n4809), .B2(
        reg_file[311]), .ZN(n6289) );
  AOI22_X1 U5944 ( .A1(n3286), .A2(reg_file[375]), .B1(n3359), .B2(
        reg_file[343]), .ZN(n6290) );
  AOI22_X1 U5945 ( .A1(n3356), .A2(reg_file[471]), .B1(n4795), .B2(
        reg_file[439]), .ZN(n6291) );
  AOI22_X1 U5946 ( .A1(n3355), .A2(reg_file[407]), .B1(n4814), .B2(
        reg_file[503]), .ZN(n6292) );
  NAND2_X1 U5947 ( .A1(n6288), .A2(n6373), .ZN(n6295) );
  NAND4_X1 U5948 ( .A1(n6287), .A2(n6286), .A3(n6285), .A4(n6284), .ZN(n6288)
         );
  AOI22_X1 U5949 ( .A1(n3358), .A2(reg_file[23]), .B1(n4809), .B2(reg_file[55]), .ZN(n6284) );
  AOI22_X1 U5950 ( .A1(n3285), .A2(reg_file[119]), .B1(n3359), .B2(
        reg_file[87]), .ZN(n6285) );
  AOI22_X1 U5951 ( .A1(n3356), .A2(reg_file[215]), .B1(n4795), .B2(
        reg_file[183]), .ZN(n6286) );
  AOI22_X1 U5952 ( .A1(n3355), .A2(reg_file[151]), .B1(n3293), .B2(
        reg_file[247]), .ZN(n6287) );
  NAND2_X1 U5953 ( .A1(n6283), .A2(n3362), .ZN(n6296) );
  NAND4_X1 U5954 ( .A1(n6282), .A2(n6281), .A3(n6280), .A4(n6279), .ZN(n6283)
         );
  AOI22_X1 U5955 ( .A1(n3358), .A2(reg_file[791]), .B1(n4808), .B2(
        reg_file[823]), .ZN(n6279) );
  AOI22_X1 U5956 ( .A1(n3285), .A2(reg_file[887]), .B1(n3359), .B2(
        reg_file[855]), .ZN(n6280) );
  AOI22_X1 U5957 ( .A1(n3356), .A2(reg_file[983]), .B1(n4795), .B2(
        reg_file[951]), .ZN(n6281) );
  AOI22_X1 U5958 ( .A1(n4790), .A2(reg_file[919]), .B1(n4815), .B2(
        reg_file[1015]), .ZN(n6282) );
  NAND2_X1 U5959 ( .A1(n6278), .A2(n3388), .ZN(n6297) );
  NAND4_X1 U5960 ( .A1(n6277), .A2(n6276), .A3(n6275), .A4(n6274), .ZN(n6278)
         );
  AOI22_X1 U5961 ( .A1(n3358), .A2(reg_file[535]), .B1(n4807), .B2(
        reg_file[567]), .ZN(n6274) );
  AOI22_X1 U5962 ( .A1(n3286), .A2(reg_file[631]), .B1(n3359), .B2(
        reg_file[599]), .ZN(n6275) );
  AOI22_X1 U5963 ( .A1(n3356), .A2(reg_file[727]), .B1(n4795), .B2(
        reg_file[695]), .ZN(n6276) );
  AOI22_X1 U5964 ( .A1(n3386), .A2(reg_file[663]), .B1(n3354), .B2(
        reg_file[759]), .ZN(n6277) );
  NAND2_X1 U5965 ( .A1(n5655), .A2(n3390), .ZN(n5656) );
  NAND4_X1 U5966 ( .A1(n5654), .A2(n5653), .A3(n5652), .A4(n5651), .ZN(n5655)
         );
  AOI22_X1 U5967 ( .A1(n4788), .A2(reg_file[535]), .B1(n4787), .B2(
        reg_file[567]), .ZN(n5651) );
  AOI22_X1 U5968 ( .A1(n4780), .A2(reg_file[631]), .B1(n4776), .B2(
        reg_file[599]), .ZN(n5652) );
  AOI22_X1 U5969 ( .A1(n3294), .A2(reg_file[695]), .B1(n3769), .B2(
        reg_file[663]), .ZN(n5653) );
  AOI22_X1 U5970 ( .A1(n4757), .A2(reg_file[727]), .B1(n4758), .B2(
        reg_file[759]), .ZN(n5654) );
  NAND2_X1 U5971 ( .A1(n5650), .A2(n3389), .ZN(n5657) );
  NAND4_X1 U5972 ( .A1(n5649), .A2(n5648), .A3(n5647), .A4(n5646), .ZN(n5650)
         );
  AOI22_X1 U5973 ( .A1(n4788), .A2(reg_file[279]), .B1(n4787), .B2(
        reg_file[311]), .ZN(n5646) );
  AOI22_X1 U5974 ( .A1(n4780), .A2(reg_file[375]), .B1(n4776), .B2(
        reg_file[343]), .ZN(n5647) );
  AOI22_X1 U5975 ( .A1(n3294), .A2(reg_file[439]), .B1(n3769), .B2(
        reg_file[407]), .ZN(n5648) );
  AOI22_X1 U5976 ( .A1(n4757), .A2(reg_file[471]), .B1(n4758), .B2(
        reg_file[503]), .ZN(n5649) );
  NAND2_X1 U5977 ( .A1(n5645), .A2(n3361), .ZN(n5658) );
  NAND4_X1 U5978 ( .A1(n5644), .A2(n5643), .A3(n5642), .A4(n5641), .ZN(n5645)
         );
  AOI22_X1 U5979 ( .A1(n4788), .A2(reg_file[791]), .B1(n4787), .B2(
        reg_file[823]), .ZN(n5641) );
  AOI22_X1 U5980 ( .A1(n4780), .A2(reg_file[887]), .B1(n4776), .B2(
        reg_file[855]), .ZN(n5642) );
  AOI22_X1 U5981 ( .A1(n3294), .A2(reg_file[951]), .B1(n3769), .B2(
        reg_file[919]), .ZN(n5643) );
  AOI22_X1 U5982 ( .A1(n4757), .A2(reg_file[983]), .B1(n4758), .B2(
        reg_file[1015]), .ZN(n5644) );
  NAND2_X1 U5983 ( .A1(n5640), .A2(n4754), .ZN(n5659) );
  NAND4_X1 U5984 ( .A1(n5639), .A2(n5638), .A3(n5637), .A4(n5636), .ZN(n5640)
         );
  AOI22_X1 U5985 ( .A1(n4788), .A2(reg_file[23]), .B1(n4786), .B2(reg_file[55]), .ZN(n5636) );
  AOI22_X1 U5986 ( .A1(n4780), .A2(reg_file[119]), .B1(n4776), .B2(
        reg_file[87]), .ZN(n5637) );
  AOI22_X1 U5987 ( .A1(n3294), .A2(reg_file[183]), .B1(n3769), .B2(
        reg_file[151]), .ZN(n5638) );
  AOI22_X1 U5988 ( .A1(n4757), .A2(reg_file[215]), .B1(n4758), .B2(
        reg_file[247]), .ZN(n5639) );
  NAND4_X1 U5989 ( .A1(n5683), .A2(n5682), .A3(n5681), .A4(n5680), .ZN(
        rs2_val_gpr_w[24]) );
  NAND2_X1 U5990 ( .A1(n5679), .A2(n4816), .ZN(n5680) );
  NAND4_X1 U5991 ( .A1(n5678), .A2(n5677), .A3(n5676), .A4(n5675), .ZN(n5679)
         );
  AOI22_X1 U5992 ( .A1(n4788), .A2(reg_file[792]), .B1(n4787), .B2(
        reg_file[824]), .ZN(n5675) );
  AOI22_X1 U5993 ( .A1(n4780), .A2(reg_file[888]), .B1(n3799), .B2(
        reg_file[856]), .ZN(n5676) );
  AOI22_X1 U5994 ( .A1(n4818), .A2(reg_file[952]), .B1(n4767), .B2(
        reg_file[920]), .ZN(n5677) );
  AOI22_X1 U5995 ( .A1(n3519), .A2(reg_file[984]), .B1(n4759), .B2(
        reg_file[1016]), .ZN(n5678) );
  NAND2_X1 U5996 ( .A1(n5674), .A2(n5804), .ZN(n5681) );
  NAND4_X1 U5997 ( .A1(n5673), .A2(n5672), .A3(n5671), .A4(n5670), .ZN(n5674)
         );
  AOI22_X1 U5998 ( .A1(n4788), .A2(reg_file[280]), .B1(n4787), .B2(
        reg_file[312]), .ZN(n5670) );
  AOI22_X1 U5999 ( .A1(n4780), .A2(reg_file[376]), .B1(n3799), .B2(
        reg_file[344]), .ZN(n5671) );
  AOI22_X1 U6000 ( .A1(n4818), .A2(reg_file[440]), .B1(n4767), .B2(
        reg_file[408]), .ZN(n5672) );
  AOI22_X1 U6001 ( .A1(n4757), .A2(reg_file[472]), .B1(n4758), .B2(
        reg_file[504]), .ZN(n5673) );
  NAND2_X1 U6002 ( .A1(n5669), .A2(n5808), .ZN(n5682) );
  NAND4_X1 U6003 ( .A1(n5668), .A2(n5667), .A3(n5666), .A4(n5665), .ZN(n5669)
         );
  AOI22_X1 U6004 ( .A1(n4788), .A2(reg_file[536]), .B1(n4786), .B2(
        reg_file[568]), .ZN(n5665) );
  AOI22_X1 U6005 ( .A1(n4780), .A2(reg_file[632]), .B1(n3799), .B2(
        reg_file[600]), .ZN(n5666) );
  AOI22_X1 U6006 ( .A1(n4818), .A2(reg_file[696]), .B1(n4767), .B2(
        reg_file[664]), .ZN(n5667) );
  AOI22_X1 U6007 ( .A1(n4757), .A2(reg_file[728]), .B1(n4759), .B2(
        reg_file[760]), .ZN(n5668) );
  NAND2_X1 U6008 ( .A1(n5664), .A2(n5805), .ZN(n5683) );
  NAND4_X1 U6009 ( .A1(n5663), .A2(n5662), .A3(n5661), .A4(n5660), .ZN(n5664)
         );
  AOI22_X1 U6010 ( .A1(n4788), .A2(reg_file[24]), .B1(n4787), .B2(reg_file[56]), .ZN(n5660) );
  AOI22_X1 U6011 ( .A1(n4780), .A2(reg_file[120]), .B1(n3799), .B2(
        reg_file[88]), .ZN(n5661) );
  AOI22_X1 U6012 ( .A1(n4818), .A2(reg_file[184]), .B1(n4767), .B2(
        reg_file[152]), .ZN(n5662) );
  AOI22_X1 U6013 ( .A1(n4757), .A2(reg_file[216]), .B1(n4759), .B2(
        reg_file[248]), .ZN(n5663) );
  AOI22_X1 U6014 ( .A1(n4812), .A2(reg_file[793]), .B1(n4809), .B2(
        reg_file[825]), .ZN(n6305) );
  AOI22_X1 U6015 ( .A1(n3286), .A2(reg_file[889]), .B1(n4805), .B2(
        reg_file[857]), .ZN(n6306) );
  AOI22_X1 U6016 ( .A1(n4800), .A2(reg_file[985]), .B1(n3360), .B2(
        reg_file[953]), .ZN(n6307) );
  AOI22_X1 U6017 ( .A1(n3355), .A2(reg_file[921]), .B1(n4814), .B2(
        reg_file[1017]), .ZN(n6308) );
  AOI22_X1 U6018 ( .A1(n4812), .A2(reg_file[537]), .B1(n4809), .B2(
        reg_file[569]), .ZN(n6301) );
  AOI22_X1 U6019 ( .A1(n3285), .A2(reg_file[633]), .B1(n4805), .B2(
        reg_file[601]), .ZN(n6302) );
  AOI22_X1 U6020 ( .A1(n4800), .A2(reg_file[729]), .B1(n3360), .B2(
        reg_file[697]), .ZN(n6303) );
  AOI22_X1 U6021 ( .A1(n3386), .A2(reg_file[665]), .B1(n4813), .B2(
        reg_file[761]), .ZN(n6304) );
  AOI22_X1 U6022 ( .A1(n3285), .A2(reg_file[377]), .B1(n4805), .B2(
        reg_file[345]), .ZN(n6298) );
  AOI22_X1 U6023 ( .A1(n4800), .A2(reg_file[473]), .B1(n3360), .B2(
        reg_file[441]), .ZN(n6299) );
  AOI22_X1 U6024 ( .A1(n3355), .A2(reg_file[409]), .B1(n3293), .B2(
        reg_file[505]), .ZN(n6300) );
  NAND4_X1 U6025 ( .A1(n6332), .A2(n6331), .A3(n6330), .A4(n6329), .ZN(
        rs1_val_gpr_w[26]) );
  NAND2_X1 U6026 ( .A1(n6328), .A2(n3388), .ZN(n6329) );
  NAND4_X1 U6027 ( .A1(n6327), .A2(n6326), .A3(n6325), .A4(n6324), .ZN(n6328)
         );
  AOI22_X1 U6028 ( .A1(n4811), .A2(reg_file[538]), .B1(n4809), .B2(
        reg_file[570]), .ZN(n6324) );
  AOI22_X1 U6029 ( .A1(n3285), .A2(reg_file[634]), .B1(n4805), .B2(
        reg_file[602]), .ZN(n6325) );
  AOI22_X1 U6030 ( .A1(n4800), .A2(reg_file[730]), .B1(n3360), .B2(
        reg_file[698]), .ZN(n6326) );
  AOI22_X1 U6031 ( .A1(n4790), .A2(reg_file[666]), .B1(n4813), .B2(
        reg_file[762]), .ZN(n6327) );
  NAND2_X1 U6032 ( .A1(n6323), .A2(n6373), .ZN(n6330) );
  NAND4_X1 U6033 ( .A1(n6322), .A2(n6321), .A3(n6320), .A4(n6319), .ZN(n6323)
         );
  AOI22_X1 U6034 ( .A1(n4812), .A2(reg_file[26]), .B1(n4809), .B2(reg_file[58]), .ZN(n6319) );
  AOI22_X1 U6035 ( .A1(n3286), .A2(reg_file[122]), .B1(n4805), .B2(
        reg_file[90]), .ZN(n6320) );
  AOI22_X1 U6036 ( .A1(n4800), .A2(reg_file[218]), .B1(n3360), .B2(
        reg_file[186]), .ZN(n6321) );
  AOI22_X1 U6037 ( .A1(n3355), .A2(reg_file[154]), .B1(n3293), .B2(
        reg_file[250]), .ZN(n6322) );
  NAND2_X1 U6038 ( .A1(n6318), .A2(n3362), .ZN(n6331) );
  NAND4_X1 U6039 ( .A1(n6317), .A2(n6316), .A3(n6315), .A4(n6314), .ZN(n6318)
         );
  AOI22_X1 U6040 ( .A1(n4812), .A2(reg_file[794]), .B1(n4809), .B2(
        reg_file[826]), .ZN(n6314) );
  AOI22_X1 U6041 ( .A1(n3286), .A2(reg_file[890]), .B1(n4805), .B2(
        reg_file[858]), .ZN(n6315) );
  AOI22_X1 U6042 ( .A1(n4800), .A2(reg_file[986]), .B1(n3360), .B2(
        reg_file[954]), .ZN(n6316) );
  AOI22_X1 U6043 ( .A1(n3355), .A2(reg_file[922]), .B1(n4814), .B2(
        reg_file[1018]), .ZN(n6317) );
  NAND2_X1 U6044 ( .A1(n6313), .A2(n3387), .ZN(n6332) );
  NAND4_X1 U6045 ( .A1(n6312), .A2(n6311), .A3(n6310), .A4(n6309), .ZN(n6313)
         );
  AOI22_X1 U6046 ( .A1(n4811), .A2(reg_file[282]), .B1(n4809), .B2(
        reg_file[314]), .ZN(n6309) );
  AOI22_X1 U6047 ( .A1(n3285), .A2(reg_file[378]), .B1(n4805), .B2(
        reg_file[346]), .ZN(n6310) );
  AOI22_X1 U6048 ( .A1(n4800), .A2(reg_file[474]), .B1(n3360), .B2(
        reg_file[442]), .ZN(n6311) );
  AOI22_X1 U6049 ( .A1(n3355), .A2(reg_file[410]), .B1(n4813), .B2(
        reg_file[506]), .ZN(n6312) );
  NAND4_X1 U6050 ( .A1(n5707), .A2(n5706), .A3(n5705), .A4(n5704), .ZN(
        rs2_val_gpr_w[26]) );
  NAND2_X1 U6051 ( .A1(n5703), .A2(n4816), .ZN(n5704) );
  NAND4_X1 U6052 ( .A1(n5702), .A2(n5701), .A3(n5700), .A4(n5699), .ZN(n5703)
         );
  AOI22_X1 U6053 ( .A1(n4788), .A2(reg_file[794]), .B1(n4787), .B2(
        reg_file[826]), .ZN(n5699) );
  AOI22_X1 U6054 ( .A1(n4779), .A2(reg_file[890]), .B1(n3799), .B2(
        reg_file[858]), .ZN(n5700) );
  AOI22_X1 U6055 ( .A1(n4818), .A2(reg_file[954]), .B1(n4767), .B2(
        reg_file[922]), .ZN(n5701) );
  AOI22_X1 U6056 ( .A1(n4757), .A2(reg_file[986]), .B1(n4759), .B2(
        reg_file[1018]), .ZN(n5702) );
  NAND2_X1 U6057 ( .A1(n5698), .A2(n5804), .ZN(n5705) );
  NAND4_X1 U6058 ( .A1(n5697), .A2(n5696), .A3(n5695), .A4(n5694), .ZN(n5698)
         );
  AOI22_X1 U6059 ( .A1(n4788), .A2(reg_file[282]), .B1(n4787), .B2(
        reg_file[314]), .ZN(n5694) );
  AOI22_X1 U6060 ( .A1(n4779), .A2(reg_file[378]), .B1(n3799), .B2(
        reg_file[346]), .ZN(n5695) );
  AOI22_X1 U6061 ( .A1(n4818), .A2(reg_file[442]), .B1(n4767), .B2(
        reg_file[410]), .ZN(n5696) );
  AOI22_X1 U6062 ( .A1(n4757), .A2(reg_file[474]), .B1(n4758), .B2(
        reg_file[506]), .ZN(n5697) );
  NAND2_X1 U6063 ( .A1(n5693), .A2(n5808), .ZN(n5706) );
  NAND4_X1 U6064 ( .A1(n5692), .A2(n5691), .A3(n5690), .A4(n5689), .ZN(n5693)
         );
  AOI22_X1 U6065 ( .A1(n4788), .A2(reg_file[538]), .B1(n4786), .B2(
        reg_file[570]), .ZN(n5689) );
  AOI22_X1 U6066 ( .A1(n4779), .A2(reg_file[634]), .B1(n3799), .B2(
        reg_file[602]), .ZN(n5690) );
  AOI22_X1 U6067 ( .A1(n4818), .A2(reg_file[698]), .B1(n4767), .B2(
        reg_file[666]), .ZN(n5691) );
  AOI22_X1 U6068 ( .A1(n4757), .A2(reg_file[730]), .B1(n4758), .B2(
        reg_file[762]), .ZN(n5692) );
  NAND2_X1 U6069 ( .A1(n5688), .A2(n5805), .ZN(n5707) );
  NAND4_X1 U6070 ( .A1(n5687), .A2(n5686), .A3(n5685), .A4(n5684), .ZN(n5688)
         );
  AOI22_X1 U6071 ( .A1(n4788), .A2(reg_file[26]), .B1(n4787), .B2(reg_file[58]), .ZN(n5684) );
  AOI22_X1 U6072 ( .A1(n4779), .A2(reg_file[122]), .B1(n3799), .B2(
        reg_file[90]), .ZN(n5685) );
  AOI22_X1 U6073 ( .A1(n4818), .A2(reg_file[186]), .B1(n4767), .B2(
        reg_file[154]), .ZN(n5686) );
  BUF_X1 U6074 ( .A(n3769), .Z(n4767) );
  AOI22_X1 U6075 ( .A1(n4755), .A2(reg_file[218]), .B1(n4759), .B2(
        reg_file[250]), .ZN(n5687) );
  AOI22_X1 U6076 ( .A1(n4801), .A2(reg_file[475]), .B1(n4796), .B2(
        reg_file[443]), .ZN(n6337) );
  AOI22_X1 U6077 ( .A1(n3386), .A2(reg_file[411]), .B1(n3293), .B2(
        reg_file[507]), .ZN(n6338) );
  AOI22_X1 U6078 ( .A1(n4811), .A2(reg_file[795]), .B1(n4809), .B2(
        reg_file[827]), .ZN(n6333) );
  AOI22_X1 U6079 ( .A1(n3286), .A2(reg_file[891]), .B1(n4806), .B2(
        reg_file[859]), .ZN(n6334) );
  AOI22_X1 U6080 ( .A1(n4801), .A2(reg_file[987]), .B1(n4796), .B2(
        reg_file[955]), .ZN(n6335) );
  AOI22_X1 U6081 ( .A1(n3355), .A2(reg_file[923]), .B1(n4813), .B2(
        reg_file[1019]), .ZN(n6336) );
  NAND4_X1 U6082 ( .A1(n5731), .A2(n5730), .A3(n5729), .A4(n5728), .ZN(
        rs2_val_gpr_w[27]) );
  NAND2_X1 U6083 ( .A1(n5727), .A2(n4816), .ZN(n5728) );
  NAND4_X1 U6084 ( .A1(n5726), .A2(n5725), .A3(n5724), .A4(n5723), .ZN(n5727)
         );
  AOI22_X1 U6085 ( .A1(n4788), .A2(reg_file[795]), .B1(n4787), .B2(
        reg_file[827]), .ZN(n5723) );
  AOI22_X1 U6086 ( .A1(n4779), .A2(reg_file[891]), .B1(n4777), .B2(
        reg_file[859]), .ZN(n5724) );
  AOI22_X1 U6087 ( .A1(n4818), .A2(reg_file[955]), .B1(n4768), .B2(
        reg_file[923]), .ZN(n5725) );
  AOI22_X1 U6088 ( .A1(n5809), .A2(reg_file[987]), .B1(n4758), .B2(
        reg_file[1019]), .ZN(n5726) );
  NAND2_X1 U6089 ( .A1(n5722), .A2(n5805), .ZN(n5729) );
  NAND4_X1 U6090 ( .A1(n5721), .A2(n5720), .A3(n5719), .A4(n5718), .ZN(n5722)
         );
  AOI22_X1 U6091 ( .A1(n4788), .A2(reg_file[27]), .B1(n4787), .B2(reg_file[59]), .ZN(n5718) );
  AOI22_X1 U6092 ( .A1(n4779), .A2(reg_file[123]), .B1(n4777), .B2(
        reg_file[91]), .ZN(n5719) );
  AOI22_X1 U6093 ( .A1(n4818), .A2(reg_file[187]), .B1(n4768), .B2(
        reg_file[155]), .ZN(n5720) );
  AOI22_X1 U6094 ( .A1(n3519), .A2(reg_file[219]), .B1(n4758), .B2(
        reg_file[251]), .ZN(n5721) );
  NAND2_X1 U6095 ( .A1(n5717), .A2(n5808), .ZN(n5730) );
  NAND4_X1 U6096 ( .A1(n5716), .A2(n5715), .A3(n5714), .A4(n5713), .ZN(n5717)
         );
  AOI22_X1 U6097 ( .A1(n4788), .A2(reg_file[539]), .B1(n4787), .B2(
        reg_file[571]), .ZN(n5713) );
  AOI22_X1 U6098 ( .A1(n4779), .A2(reg_file[635]), .B1(n4777), .B2(
        reg_file[603]), .ZN(n5714) );
  AOI22_X1 U6099 ( .A1(n4818), .A2(reg_file[699]), .B1(n4768), .B2(
        reg_file[667]), .ZN(n5715) );
  AOI22_X1 U6100 ( .A1(n4757), .A2(reg_file[731]), .B1(n4758), .B2(
        reg_file[763]), .ZN(n5716) );
  NAND2_X1 U6101 ( .A1(n5712), .A2(n5804), .ZN(n5731) );
  NAND4_X1 U6102 ( .A1(n5711), .A2(n5710), .A3(n5709), .A4(n5708), .ZN(n5712)
         );
  AOI22_X1 U6103 ( .A1(n4788), .A2(reg_file[283]), .B1(n4786), .B2(
        reg_file[315]), .ZN(n5708) );
  AOI22_X1 U6104 ( .A1(n4779), .A2(reg_file[379]), .B1(n4777), .B2(
        reg_file[347]), .ZN(n5709) );
  AOI22_X1 U6105 ( .A1(n4818), .A2(reg_file[443]), .B1(n4768), .B2(
        reg_file[411]), .ZN(n5710) );
  AOI22_X1 U6106 ( .A1(n4756), .A2(reg_file[475]), .B1(n4758), .B2(
        reg_file[507]), .ZN(n5711) );
  NAND4_X1 U6107 ( .A1(n5755), .A2(n5754), .A3(n5753), .A4(n5752), .ZN(
        rs2_val_gpr_w[28]) );
  NAND2_X1 U6108 ( .A1(n5751), .A2(n5808), .ZN(n5752) );
  NAND4_X1 U6109 ( .A1(n5750), .A2(n5749), .A3(n5748), .A4(n5747), .ZN(n5751)
         );
  AOI22_X1 U6110 ( .A1(n4788), .A2(reg_file[540]), .B1(n4787), .B2(
        reg_file[572]), .ZN(n5747) );
  AOI22_X1 U6111 ( .A1(n4778), .A2(reg_file[636]), .B1(n4777), .B2(
        reg_file[604]), .ZN(n5748) );
  AOI22_X1 U6112 ( .A1(n4818), .A2(reg_file[700]), .B1(n4768), .B2(
        reg_file[668]), .ZN(n5749) );
  AOI22_X1 U6113 ( .A1(n4757), .A2(reg_file[732]), .B1(n4758), .B2(
        reg_file[764]), .ZN(n5750) );
  NAND2_X1 U6114 ( .A1(n5746), .A2(n5805), .ZN(n5753) );
  NAND4_X1 U6115 ( .A1(n5745), .A2(n5744), .A3(n5743), .A4(n5742), .ZN(n5746)
         );
  AOI22_X1 U6116 ( .A1(n4788), .A2(reg_file[28]), .B1(n4787), .B2(reg_file[60]), .ZN(n5742) );
  AOI22_X1 U6117 ( .A1(n4779), .A2(reg_file[124]), .B1(n4777), .B2(
        reg_file[92]), .ZN(n5743) );
  AOI22_X1 U6118 ( .A1(n4818), .A2(reg_file[188]), .B1(n4768), .B2(
        reg_file[156]), .ZN(n5744) );
  AOI22_X1 U6119 ( .A1(n4757), .A2(reg_file[220]), .B1(n4758), .B2(
        reg_file[252]), .ZN(n5745) );
  NAND2_X1 U6120 ( .A1(n5741), .A2(n4816), .ZN(n5754) );
  NAND4_X1 U6121 ( .A1(n5740), .A2(n5739), .A3(n5738), .A4(n5737), .ZN(n5741)
         );
  AOI22_X1 U6122 ( .A1(n4788), .A2(reg_file[796]), .B1(n4787), .B2(
        reg_file[828]), .ZN(n5737) );
  AOI22_X1 U6123 ( .A1(n4779), .A2(reg_file[892]), .B1(n4777), .B2(
        reg_file[860]), .ZN(n5738) );
  AOI22_X1 U6124 ( .A1(n4818), .A2(reg_file[956]), .B1(n4768), .B2(
        reg_file[924]), .ZN(n5739) );
  AOI22_X1 U6125 ( .A1(n4757), .A2(reg_file[988]), .B1(n4758), .B2(
        reg_file[1020]), .ZN(n5740) );
  NAND2_X1 U6126 ( .A1(n5736), .A2(n5804), .ZN(n5755) );
  NAND4_X1 U6127 ( .A1(n5735), .A2(n5734), .A3(n5733), .A4(n5732), .ZN(n5736)
         );
  AOI22_X1 U6128 ( .A1(n4788), .A2(reg_file[284]), .B1(n4787), .B2(
        reg_file[316]), .ZN(n5732) );
  AOI22_X1 U6129 ( .A1(n4779), .A2(reg_file[380]), .B1(n4777), .B2(
        reg_file[348]), .ZN(n5733) );
  AOI22_X1 U6130 ( .A1(n4818), .A2(reg_file[444]), .B1(n4768), .B2(
        reg_file[412]), .ZN(n5734) );
  AOI22_X1 U6131 ( .A1(n5809), .A2(reg_file[476]), .B1(n4758), .B2(
        reg_file[508]), .ZN(n5735) );
  NAND2_X1 U6132 ( .A1(n6358), .A2(n3362), .ZN(n6359) );
  NAND4_X1 U6133 ( .A1(n6357), .A2(n6356), .A3(n6355), .A4(n6354), .ZN(n6358)
         );
  AOI22_X1 U6134 ( .A1(n4812), .A2(reg_file[797]), .B1(n4809), .B2(
        reg_file[829]), .ZN(n6354) );
  AOI22_X1 U6135 ( .A1(n3285), .A2(reg_file[893]), .B1(n4806), .B2(
        reg_file[861]), .ZN(n6355) );
  AOI22_X1 U6136 ( .A1(n4801), .A2(reg_file[989]), .B1(n4796), .B2(
        reg_file[957]), .ZN(n6356) );
  AOI22_X1 U6137 ( .A1(reg_file[925]), .A2(n3355), .B1(n4814), .B2(
        reg_file[1021]), .ZN(n6357) );
  NAND2_X1 U6138 ( .A1(n6353), .A2(n6373), .ZN(n6360) );
  NAND4_X1 U6139 ( .A1(n6352), .A2(n6351), .A3(n6350), .A4(n6349), .ZN(n6353)
         );
  AOI22_X1 U6140 ( .A1(n4811), .A2(reg_file[29]), .B1(n4809), .B2(reg_file[61]), .ZN(n6349) );
  AOI22_X1 U6141 ( .A1(n3285), .A2(reg_file[125]), .B1(n4806), .B2(
        reg_file[93]), .ZN(n6350) );
  AOI22_X1 U6142 ( .A1(n4801), .A2(reg_file[221]), .B1(n4796), .B2(
        reg_file[189]), .ZN(n6351) );
  AOI22_X1 U6143 ( .A1(n3386), .A2(reg_file[157]), .B1(n4813), .B2(
        reg_file[253]), .ZN(n6352) );
  NAND2_X1 U6144 ( .A1(n6348), .A2(n3387), .ZN(n6361) );
  NAND4_X1 U6145 ( .A1(n6347), .A2(n6346), .A3(n6345), .A4(n6344), .ZN(n6348)
         );
  AOI22_X1 U6146 ( .A1(n4812), .A2(reg_file[285]), .B1(n4809), .B2(
        reg_file[317]), .ZN(n6344) );
  AOI22_X1 U6147 ( .A1(n3285), .A2(reg_file[381]), .B1(n4805), .B2(
        reg_file[349]), .ZN(n6345) );
  AOI22_X1 U6148 ( .A1(n4800), .A2(reg_file[477]), .B1(n4796), .B2(
        reg_file[445]), .ZN(n6346) );
  AOI22_X1 U6149 ( .A1(n3355), .A2(reg_file[413]), .B1(n3293), .B2(
        reg_file[509]), .ZN(n6347) );
  NAND2_X1 U6150 ( .A1(n6343), .A2(n3388), .ZN(n6362) );
  NAND4_X1 U6151 ( .A1(n6342), .A2(n6341), .A3(n6340), .A4(n6339), .ZN(n6343)
         );
  AOI22_X1 U6152 ( .A1(n4811), .A2(reg_file[541]), .B1(n4809), .B2(
        reg_file[573]), .ZN(n6339) );
  AOI22_X1 U6153 ( .A1(n3286), .A2(reg_file[637]), .B1(n4805), .B2(
        reg_file[605]), .ZN(n6340) );
  AOI22_X1 U6154 ( .A1(n4800), .A2(reg_file[733]), .B1(n4796), .B2(
        reg_file[701]), .ZN(n6341) );
  AOI22_X1 U6155 ( .A1(n3355), .A2(reg_file[669]), .B1(n4814), .B2(
        reg_file[765]), .ZN(n6342) );
  NAND4_X1 U6156 ( .A1(n5779), .A2(n5778), .A3(n5777), .A4(n5776), .ZN(
        rs2_val_gpr_w[29]) );
  NAND2_X1 U6157 ( .A1(n5775), .A2(n4816), .ZN(n5776) );
  NAND4_X1 U6158 ( .A1(n5774), .A2(n5773), .A3(n5772), .A4(n5771), .ZN(n5775)
         );
  AOI22_X1 U6159 ( .A1(n4788), .A2(reg_file[797]), .B1(n4787), .B2(
        reg_file[829]), .ZN(n5771) );
  AOI22_X1 U6160 ( .A1(n4778), .A2(reg_file[893]), .B1(n4777), .B2(
        reg_file[861]), .ZN(n5772) );
  AOI22_X1 U6161 ( .A1(n4818), .A2(reg_file[957]), .B1(n4768), .B2(
        reg_file[925]), .ZN(n5773) );
  AOI22_X1 U6162 ( .A1(n4757), .A2(reg_file[989]), .B1(n4758), .B2(
        reg_file[1021]), .ZN(n5774) );
  NAND2_X1 U6163 ( .A1(n5770), .A2(n5804), .ZN(n5777) );
  NAND4_X1 U6164 ( .A1(n5769), .A2(n5768), .A3(n5767), .A4(n5766), .ZN(n5770)
         );
  AOI22_X1 U6165 ( .A1(n4788), .A2(reg_file[285]), .B1(n4787), .B2(
        reg_file[317]), .ZN(n5766) );
  AOI22_X1 U6166 ( .A1(n4778), .A2(reg_file[381]), .B1(n4777), .B2(
        reg_file[349]), .ZN(n5767) );
  AOI22_X1 U6167 ( .A1(n4818), .A2(reg_file[445]), .B1(n4768), .B2(
        reg_file[413]), .ZN(n5768) );
  AOI22_X1 U6168 ( .A1(n4756), .A2(reg_file[477]), .B1(n4758), .B2(
        reg_file[509]), .ZN(n5769) );
  NAND2_X1 U6169 ( .A1(n5765), .A2(n5808), .ZN(n5778) );
  NAND4_X1 U6170 ( .A1(n5764), .A2(n5763), .A3(n5762), .A4(n5761), .ZN(n5765)
         );
  AOI22_X1 U6171 ( .A1(n4788), .A2(reg_file[541]), .B1(n4787), .B2(
        reg_file[573]), .ZN(n5761) );
  AOI22_X1 U6172 ( .A1(n4778), .A2(reg_file[637]), .B1(n4777), .B2(
        reg_file[605]), .ZN(n5762) );
  AOI22_X1 U6173 ( .A1(n4818), .A2(reg_file[701]), .B1(n4768), .B2(
        reg_file[669]), .ZN(n5763) );
  AOI22_X1 U6174 ( .A1(n4756), .A2(reg_file[733]), .B1(n4758), .B2(
        reg_file[765]), .ZN(n5764) );
  NAND2_X1 U6175 ( .A1(n5760), .A2(n5805), .ZN(n5779) );
  NAND4_X1 U6176 ( .A1(n5759), .A2(n5758), .A3(n5757), .A4(n5756), .ZN(n5760)
         );
  AOI22_X1 U6177 ( .A1(n4788), .A2(reg_file[29]), .B1(n4787), .B2(reg_file[61]), .ZN(n5756) );
  AOI22_X1 U6178 ( .A1(n4778), .A2(reg_file[125]), .B1(n4777), .B2(
        reg_file[93]), .ZN(n5757) );
  AOI22_X1 U6179 ( .A1(n4818), .A2(reg_file[189]), .B1(n4768), .B2(
        reg_file[157]), .ZN(n5758) );
  AOI22_X1 U6180 ( .A1(n4757), .A2(reg_file[221]), .B1(n4758), .B2(
        reg_file[253]), .ZN(n5759) );
  AOI22_X1 U6181 ( .A1(n4811), .A2(reg_file[798]), .B1(n4809), .B2(
        reg_file[830]), .ZN(n6365) );
  AOI22_X1 U6182 ( .A1(n3286), .A2(reg_file[894]), .B1(n4806), .B2(
        reg_file[862]), .ZN(n6366) );
  AOI22_X1 U6183 ( .A1(n4801), .A2(reg_file[990]), .B1(n4797), .B2(
        reg_file[958]), .ZN(n6367) );
  AOI22_X1 U6184 ( .A1(n3355), .A2(reg_file[926]), .B1(n4813), .B2(
        reg_file[1022]), .ZN(n6368) );
  AOI22_X1 U6185 ( .A1(n4801), .A2(reg_file[222]), .B1(n4797), .B2(
        reg_file[190]), .ZN(n6363) );
  AOI22_X1 U6186 ( .A1(n3355), .A2(reg_file[158]), .B1(n4813), .B2(
        reg_file[254]), .ZN(n6364) );
  NAND4_X1 U6187 ( .A1(n5803), .A2(n5802), .A3(n5801), .A4(n5800), .ZN(
        rs2_val_gpr_w[30]) );
  NAND2_X1 U6188 ( .A1(n5799), .A2(n4816), .ZN(n5800) );
  NAND4_X1 U6189 ( .A1(n5798), .A2(n5797), .A3(n5796), .A4(n5795), .ZN(n5799)
         );
  AOI22_X1 U6190 ( .A1(n4788), .A2(reg_file[798]), .B1(n4787), .B2(
        reg_file[830]), .ZN(n5795) );
  AOI22_X1 U6191 ( .A1(n4778), .A2(reg_file[894]), .B1(n3799), .B2(
        reg_file[862]), .ZN(n5796) );
  AOI22_X1 U6192 ( .A1(n4818), .A2(reg_file[958]), .B1(n3769), .B2(
        reg_file[926]), .ZN(n5797) );
  AOI22_X1 U6193 ( .A1(n4757), .A2(reg_file[990]), .B1(n4758), .B2(
        reg_file[1022]), .ZN(n5798) );
  NAND2_X1 U6194 ( .A1(n5794), .A2(n5804), .ZN(n5801) );
  NAND4_X1 U6195 ( .A1(n5793), .A2(n5792), .A3(n5791), .A4(n5790), .ZN(n5794)
         );
  AOI22_X1 U6196 ( .A1(n4788), .A2(reg_file[286]), .B1(n4787), .B2(
        reg_file[318]), .ZN(n5790) );
  AOI22_X1 U6197 ( .A1(n4778), .A2(reg_file[382]), .B1(n3799), .B2(
        reg_file[350]), .ZN(n5791) );
  AOI22_X1 U6198 ( .A1(n4818), .A2(reg_file[446]), .B1(n3769), .B2(
        reg_file[414]), .ZN(n5792) );
  AOI22_X1 U6199 ( .A1(n4756), .A2(reg_file[478]), .B1(n4758), .B2(
        reg_file[510]), .ZN(n5793) );
  NAND2_X1 U6200 ( .A1(n5789), .A2(n5808), .ZN(n5802) );
  NAND4_X1 U6201 ( .A1(n5788), .A2(n5787), .A3(n5786), .A4(n5785), .ZN(n5789)
         );
  AOI22_X1 U6202 ( .A1(n4788), .A2(reg_file[542]), .B1(n4787), .B2(
        reg_file[574]), .ZN(n5785) );
  AOI22_X1 U6203 ( .A1(n4778), .A2(reg_file[638]), .B1(n3799), .B2(
        reg_file[606]), .ZN(n5786) );
  AOI22_X1 U6204 ( .A1(n4818), .A2(reg_file[702]), .B1(n3769), .B2(
        reg_file[670]), .ZN(n5787) );
  AOI22_X1 U6205 ( .A1(n4756), .A2(reg_file[734]), .B1(n4758), .B2(
        reg_file[766]), .ZN(n5788) );
  NAND2_X1 U6206 ( .A1(n5784), .A2(n5805), .ZN(n5803) );
  NAND4_X1 U6207 ( .A1(n5783), .A2(n5782), .A3(n5781), .A4(n5780), .ZN(n5784)
         );
  AOI22_X1 U6208 ( .A1(n4788), .A2(reg_file[30]), .B1(n4787), .B2(reg_file[62]), .ZN(n5780) );
  NOR2_X1 U6209 ( .A1(n4976), .A2(n6623), .ZN(n5813) );
  NAND2_X1 U6210 ( .A1(mem_i_inst_i[21]), .A2(mem_i_inst_i[22]), .ZN(n4976) );
  AOI22_X1 U6211 ( .A1(n4778), .A2(reg_file[126]), .B1(n3799), .B2(
        reg_file[94]), .ZN(n5781) );
  NOR2_X1 U6212 ( .A1(mem_i_inst_i[21]), .A2(mem_i_inst_i[20]), .ZN(n4975) );
  AOI22_X1 U6213 ( .A1(n4818), .A2(reg_file[190]), .B1(n3769), .B2(
        reg_file[158]), .ZN(n5782) );
  INV_X1 U6214 ( .A(mem_i_inst_i[22]), .ZN(n6410) );
  AOI22_X1 U6215 ( .A1(n4755), .A2(reg_file[222]), .B1(n4759), .B2(
        reg_file[254]), .ZN(n5783) );
  XNOR2_X1 U6216 ( .A(n6393), .B(n6474), .ZN(n6770) );
  INV_X1 U6217 ( .A(reset_vector_i[31]), .ZN(n6474) );
  NAND2_X1 U6218 ( .A1(n6481), .A2(reset_vector_i[30]), .ZN(n6393) );
  NOR2_X1 U6219 ( .A1(n6482), .A2(n6483), .ZN(n6481) );
  INV_X1 U6220 ( .A(reset_vector_i[29]), .ZN(n6483) );
  NAND2_X1 U6221 ( .A1(n6494), .A2(reset_vector_i[28]), .ZN(n6482) );
  NOR2_X1 U6222 ( .A1(n6496), .A2(n6495), .ZN(n6494) );
  INV_X1 U6223 ( .A(reset_vector_i[27]), .ZN(n6495) );
  NAND2_X1 U6224 ( .A1(n6507), .A2(reset_vector_i[26]), .ZN(n6496) );
  NOR2_X1 U6225 ( .A1(n6687), .A2(n6505), .ZN(n6507) );
  INV_X1 U6226 ( .A(reset_vector_i[25]), .ZN(n6505) );
  NAND2_X1 U6227 ( .A1(n6870), .A2(n6473), .ZN(n6468) );
  INV_X1 U6228 ( .A(n6760), .ZN(n6473) );
  INV_X1 U6229 ( .A(n6460), .ZN(n6472) );
  NOR2_X1 U6230 ( .A1(exception_w), .A2(n6415), .ZN(n6460) );
  AOI211_X1 U6231 ( .C1(n6757), .C2(n6844), .A(n6759), .B(n6672), .ZN(n6674)
         );
  NOR2_X1 U6232 ( .A1(n6854), .A2(n7990), .ZN(n6672) );
  NAND2_X1 U6233 ( .A1(n6395), .A2(mem_i_inst_i[12]), .ZN(n6854) );
  INV_X1 U6234 ( .A(n6873), .ZN(n6395) );
  INV_X1 U6235 ( .A(n6759), .ZN(n6675) );
  AOI22_X1 U6236 ( .A1(n7990), .A2(n6623), .B1(n7986), .B2(n7992), .ZN(
        u_lsu_N14) );
  NAND4_X1 U6237 ( .A1(n4964), .A2(n4963), .A3(n4962), .A4(n4961), .ZN(n4965)
         );
  NAND2_X1 U6238 ( .A1(n4960), .A2(n6392), .ZN(n4967) );
  NAND4_X1 U6239 ( .A1(n4959), .A2(n4958), .A3(n4957), .A4(n4956), .ZN(n4960)
         );
  NAND2_X1 U6240 ( .A1(n4955), .A2(n3362), .ZN(n4968) );
  NAND4_X1 U6241 ( .A1(n4954), .A2(n4953), .A3(n4952), .A4(n4951), .ZN(n4955)
         );
  NAND2_X1 U6242 ( .A1(n4950), .A2(n6373), .ZN(n4969) );
  NAND4_X1 U6243 ( .A1(n4949), .A2(n4948), .A3(n4947), .A4(n4946), .ZN(n4950)
         );
  AOI22_X1 U6244 ( .A1(n7990), .A2(n6411), .B1(n7988), .B2(n7992), .ZN(
        add_x_67_B_1_) );
  INV_X1 U6245 ( .A(mem_i_inst_i[21]), .ZN(n6411) );
  NAND2_X1 U6246 ( .A1(n5837), .A2(n6381), .ZN(n5838) );
  NAND4_X1 U6247 ( .A1(n5836), .A2(n5835), .A3(n5834), .A4(n5833), .ZN(n5837)
         );
  NAND2_X1 U6248 ( .A1(n5832), .A2(n6373), .ZN(n5839) );
  NAND4_X1 U6249 ( .A1(n5831), .A2(n5830), .A3(n5829), .A4(n5828), .ZN(n5832)
         );
  NAND2_X1 U6250 ( .A1(n5827), .A2(n3362), .ZN(n5840) );
  NAND4_X1 U6251 ( .A1(n5826), .A2(n5825), .A3(n5824), .A4(n5823), .ZN(n5827)
         );
  NAND2_X1 U6252 ( .A1(n5822), .A2(n6392), .ZN(n5841) );
  NAND4_X1 U6253 ( .A1(n5821), .A2(n5820), .A3(n5819), .A4(n5818), .ZN(n5822)
         );
  NAND2_X1 U6254 ( .A1(mem_i_inst_i[15]), .A2(mem_i_inst_i[17]), .ZN(n4944) );
  OAI211_X1 U6255 ( .C1(mem_i_inst_i[4]), .C2(n6752), .A(n6408), .B(n6469), 
        .ZN(n6753) );
  NAND2_X1 U6256 ( .A1(n6407), .A2(n6406), .ZN(n6469) );
  NOR3_X1 U6257 ( .A1(n4817), .A2(n6567), .A3(n6405), .ZN(n6406) );
  NAND4_X1 U6258 ( .A1(mem_i_inst_i[29]), .A2(n6830), .A3(n4910), .A4(n6827), 
        .ZN(n6405) );
  INV_X1 U6259 ( .A(mem_i_inst_i[28]), .ZN(n6567) );
  NOR2_X1 U6260 ( .A1(mem_i_inst_i[22]), .A2(mem_i_inst_i[20]), .ZN(n4974) );
  INV_X1 U6261 ( .A(n6403), .ZN(n6407) );
  INV_X1 U6262 ( .A(n6415), .ZN(n6408) );
  AND2_X1 U6263 ( .A1(n6402), .A2(n6729), .ZN(n6415) );
  NOR2_X1 U6264 ( .A1(n6403), .A2(n6401), .ZN(n6402) );
  INV_X1 U6265 ( .A(n6400), .ZN(n6401) );
  NAND3_X1 U6266 ( .A1(n6728), .A2(n6681), .A3(n6399), .ZN(n6403) );
  NOR3_X1 U6267 ( .A1(n3317), .A2(n6398), .A3(n3800), .ZN(n6399) );
  NAND3_X1 U6268 ( .A1(n3362), .A2(n6564), .A3(n6824), .ZN(n6398) );
  INV_X1 U6269 ( .A(mem_i_inst_i[30]), .ZN(n6564) );
  NOR2_X1 U6270 ( .A1(mem_i_inst_i[15]), .A2(mem_i_inst_i[17]), .ZN(n4943) );
  NOR2_X1 U6271 ( .A1(n6873), .A2(mem_i_inst_i[12]), .ZN(n6681) );
  INV_X1 U6272 ( .A(mem_i_inst_i[5]), .ZN(n6748) );
  INV_X1 U6273 ( .A(n6782), .ZN(n6791) );
  NOR2_X1 U6274 ( .A1(n6457), .A2(n6747), .ZN(n6679) );
  NAND3_X1 U6275 ( .A1(n6755), .A2(mem_i_inst_i[5]), .A3(mem_i_inst_i[6]), 
        .ZN(n6457) );
  INV_X1 U6276 ( .A(n6463), .ZN(n6464) );
  AND2_X1 U6277 ( .A1(n7212), .A2(n7676), .ZN(n3864) );
  NAND2_X1 U6278 ( .A1(n4718), .A2(n6454), .ZN(n4709) );
  NAND2_X1 U6279 ( .A1(n4711), .A2(n6742), .ZN(n4710) );
  INV_X1 U6280 ( .A(n4719), .ZN(n4711) );
  NAND2_X1 U6281 ( .A1(n6453), .A2(n6452), .ZN(n4719) );
  MUX2_X1 U6314 ( .A(n3864), .B(n4752), .S(alu_a_q[9]), .Z(n7223) );
  AOI22_X1 U6315 ( .A1(n3286), .A2(reg_file[354]), .B1(n4802), .B2(
        reg_file[322]), .ZN(n5843) );
  AOI22_X1 U6316 ( .A1(n3285), .A2(reg_file[866]), .B1(n4802), .B2(
        reg_file[834]), .ZN(n5848) );
  AOI22_X1 U6317 ( .A1(n3285), .A2(reg_file[98]), .B1(n4802), .B2(reg_file[66]), .ZN(n5853) );
  AOI22_X1 U6318 ( .A1(n3286), .A2(reg_file[610]), .B1(n4802), .B2(
        reg_file[578]), .ZN(n5858) );
  AOI22_X1 U6319 ( .A1(n3286), .A2(reg_file[609]), .B1(n4802), .B2(
        reg_file[577]), .ZN(n5819) );
  AOI22_X1 U6320 ( .A1(n3285), .A2(reg_file[865]), .B1(n4802), .B2(
        reg_file[833]), .ZN(n5824) );
  AOI22_X1 U6321 ( .A1(n3285), .A2(reg_file[97]), .B1(n4802), .B2(reg_file[65]), .ZN(n5829) );
  AOI22_X1 U6322 ( .A1(n3286), .A2(reg_file[353]), .B1(n4802), .B2(
        reg_file[321]), .ZN(n5834) );
  AOI22_X1 U6323 ( .A1(n3286), .A2(reg_file[96]), .B1(n4802), .B2(reg_file[64]), .ZN(n4947) );
  AOI22_X1 U6324 ( .A1(n3285), .A2(reg_file[352]), .B1(n4802), .B2(
        reg_file[320]), .ZN(n4962) );
  AOI22_X1 U6325 ( .A1(n3285), .A2(reg_file[864]), .B1(n4802), .B2(
        reg_file[832]), .ZN(n4952) );
  AOI22_X1 U6326 ( .A1(n3286), .A2(reg_file[608]), .B1(n4802), .B2(
        reg_file[576]), .ZN(n4957) );
  AOI22_X1 U6327 ( .A1(n5811), .A2(reg_file[98]), .B1(n4769), .B2(reg_file[66]), .ZN(n5092) );
  AOI22_X1 U6328 ( .A1(n5811), .A2(reg_file[610]), .B1(n4769), .B2(
        reg_file[578]), .ZN(n5097) );
  AOI22_X1 U6329 ( .A1(n5811), .A2(reg_file[354]), .B1(n4769), .B2(
        reg_file[322]), .ZN(n5102) );
  AOI22_X1 U6330 ( .A1(n4785), .A2(reg_file[866]), .B1(n4769), .B2(
        reg_file[834]), .ZN(n5107) );
  AOI22_X1 U6331 ( .A1(n5811), .A2(reg_file[352]), .B1(n4769), .B2(
        reg_file[320]), .ZN(n4978) );
  AOI22_X1 U6332 ( .A1(n5811), .A2(reg_file[608]), .B1(n4769), .B2(
        reg_file[576]), .ZN(n4983) );
  AOI22_X1 U6333 ( .A1(n5811), .A2(reg_file[96]), .B1(n4769), .B2(reg_file[64]), .ZN(n4988) );
  AOI22_X1 U6334 ( .A1(n5811), .A2(reg_file[864]), .B1(n4769), .B2(
        reg_file[832]), .ZN(n4993) );
  AOI22_X1 U6335 ( .A1(n5811), .A2(reg_file[97]), .B1(n4769), .B2(reg_file[65]), .ZN(n5035) );
  AOI22_X1 U6336 ( .A1(n5811), .A2(reg_file[865]), .B1(n4769), .B2(
        reg_file[833]), .ZN(n5040) );
  AOI22_X1 U6337 ( .A1(n5811), .A2(reg_file[353]), .B1(n4769), .B2(
        reg_file[321]), .ZN(n5045) );
  AOI22_X1 U6338 ( .A1(n5811), .A2(reg_file[609]), .B1(n4769), .B2(
        reg_file[577]), .ZN(n5050) );
  AOI22_X1 U6339 ( .A1(n4810), .A2(reg_file[258]), .B1(n4807), .B2(
        reg_file[290]), .ZN(n5842) );
  AOI22_X1 U6340 ( .A1(n4810), .A2(reg_file[770]), .B1(n4807), .B2(
        reg_file[802]), .ZN(n5847) );
  AOI22_X1 U6341 ( .A1(n4810), .A2(reg_file[2]), .B1(n4808), .B2(reg_file[34]), 
        .ZN(n5852) );
  AOI22_X1 U6342 ( .A1(n4810), .A2(reg_file[514]), .B1(n4809), .B2(
        reg_file[546]), .ZN(n5857) );
  AOI22_X1 U6343 ( .A1(n4810), .A2(reg_file[513]), .B1(n4808), .B2(
        reg_file[545]), .ZN(n5818) );
  AOI22_X1 U6344 ( .A1(n4810), .A2(reg_file[769]), .B1(n4807), .B2(
        reg_file[801]), .ZN(n5823) );
  AOI22_X1 U6345 ( .A1(n4810), .A2(reg_file[1]), .B1(n4807), .B2(reg_file[33]), 
        .ZN(n5828) );
  AOI22_X1 U6346 ( .A1(n4810), .A2(reg_file[257]), .B1(n4808), .B2(
        reg_file[289]), .ZN(n5833) );
  AOI22_X1 U6347 ( .A1(n4810), .A2(reg_file[0]), .B1(n4809), .B2(reg_file[32]), 
        .ZN(n4946) );
  AOI22_X1 U6348 ( .A1(n4810), .A2(reg_file[256]), .B1(n4807), .B2(
        reg_file[288]), .ZN(n4961) );
  AOI22_X1 U6349 ( .A1(n4810), .A2(reg_file[768]), .B1(n4809), .B2(
        reg_file[800]), .ZN(n4951) );
  AOI22_X1 U6350 ( .A1(n4810), .A2(reg_file[512]), .B1(n4808), .B2(
        reg_file[544]), .ZN(n4956) );
  AOI22_X1 U6351 ( .A1(n6868), .A2(rs2_val_gpr_w[0]), .B1(n4822), .B2(
        mem_d_data_wr_o[0]), .ZN(n1380) );
  XNOR2_X1 U6352 ( .A(rs2_val_gpr_w[0]), .B(n3521), .ZN(n6425) );
  AOI22_X1 U6353 ( .A1(n3296), .A2(reg_file[2]), .B1(n4787), .B2(reg_file[34]), 
        .ZN(n5091) );
  AOI22_X1 U6354 ( .A1(n3296), .A2(reg_file[514]), .B1(n4787), .B2(
        reg_file[546]), .ZN(n5096) );
  AOI22_X1 U6355 ( .A1(n3296), .A2(reg_file[1]), .B1(n4787), .B2(reg_file[33]), 
        .ZN(n5034) );
  AOI22_X1 U6356 ( .A1(n3296), .A2(reg_file[258]), .B1(n4787), .B2(
        reg_file[290]), .ZN(n5101) );
  AOI22_X1 U6357 ( .A1(n3296), .A2(reg_file[770]), .B1(n4787), .B2(
        reg_file[802]), .ZN(n5106) );
  AOI22_X1 U6358 ( .A1(n3296), .A2(reg_file[769]), .B1(n4787), .B2(
        reg_file[801]), .ZN(n5039) );
  AOI22_X1 U6359 ( .A1(n3296), .A2(reg_file[257]), .B1(n4786), .B2(
        reg_file[289]), .ZN(n5044) );
  AOI22_X1 U6360 ( .A1(n3296), .A2(reg_file[513]), .B1(n4786), .B2(
        reg_file[545]), .ZN(n5049) );
  AOI22_X1 U6361 ( .A1(n3296), .A2(reg_file[256]), .B1(n4787), .B2(
        reg_file[288]), .ZN(n4977) );
  AOI22_X1 U6362 ( .A1(n3296), .A2(reg_file[512]), .B1(n4787), .B2(
        reg_file[544]), .ZN(n4982) );
  AOI22_X1 U6363 ( .A1(n3296), .A2(reg_file[0]), .B1(n4786), .B2(reg_file[32]), 
        .ZN(n4987) );
  AOI22_X1 U6364 ( .A1(n3296), .A2(reg_file[768]), .B1(n4786), .B2(
        reg_file[800]), .ZN(n4992) );
  NAND3_X1 U6365 ( .A1(U4_RSOP_173_C3_DATA1_0), .A2(n6587), .A3(n4820), .ZN(
        n6591) );
  AOI211_X1 U6366 ( .C1(n7007), .C2(rs1_val_gpr_w[2]), .A(n6594), .B(n6897), 
        .ZN(n6595) );
  XNOR2_X1 U6367 ( .A(rs2_val_gpr_w[2]), .B(rs1_val_gpr_w[2]), .ZN(n6433) );
  AOI22_X1 U6368 ( .A1(n3386), .A2(reg_file[641]), .B1(n3522), .B2(
        reg_file[737]), .ZN(n5821) );
  AOI22_X1 U6369 ( .A1(n3386), .A2(reg_file[897]), .B1(n3522), .B2(
        reg_file[993]), .ZN(n5826) );
  AOI22_X1 U6370 ( .A1(n3386), .A2(reg_file[129]), .B1(n3522), .B2(
        reg_file[225]), .ZN(n5831) );
  AOI22_X1 U6371 ( .A1(n3386), .A2(reg_file[385]), .B1(n3522), .B2(
        reg_file[481]), .ZN(n5836) );
  AOI22_X1 U6372 ( .A1(n3355), .A2(reg_file[386]), .B1(n3522), .B2(
        reg_file[482]), .ZN(n5845) );
  AOI22_X1 U6373 ( .A1(reg_file[128]), .A2(n3386), .B1(n3293), .B2(
        reg_file[224]), .ZN(n4949) );
  AOI22_X1 U6374 ( .A1(n3355), .A2(reg_file[898]), .B1(n3354), .B2(
        reg_file[994]), .ZN(n5850) );
  AOI22_X1 U6375 ( .A1(n3386), .A2(reg_file[130]), .B1(n3354), .B2(
        reg_file[226]), .ZN(n5855) );
  AOI22_X1 U6376 ( .A1(n3386), .A2(reg_file[384]), .B1(n3354), .B2(
        reg_file[480]), .ZN(n4964) );
  AOI22_X1 U6377 ( .A1(n3386), .A2(reg_file[896]), .B1(n4814), .B2(
        reg_file[992]), .ZN(n4954) );
  AOI22_X1 U6378 ( .A1(n3386), .A2(reg_file[642]), .B1(n3354), .B2(
        reg_file[738]), .ZN(n5860) );
  AOI22_X1 U6379 ( .A1(n4790), .A2(reg_file[640]), .B1(n3354), .B2(
        reg_file[736]), .ZN(n4959) );
  AOI22_X1 U6380 ( .A1(n6868), .A2(rs2_val_gpr_w[1]), .B1(n4822), .B2(
        mem_d_data_wr_o[1]), .ZN(n1381) );
  AOI22_X1 U6381 ( .A1(n3357), .A2(reg_file[162]), .B1(n4761), .B2(
        reg_file[130]), .ZN(n5093) );
  AOI22_X1 U6382 ( .A1(n3357), .A2(reg_file[416]), .B1(n4761), .B2(
        reg_file[384]), .ZN(n4979) );
  AOI22_X1 U6383 ( .A1(n3357), .A2(reg_file[674]), .B1(n4761), .B2(
        reg_file[642]), .ZN(n5098) );
  AOI22_X1 U6384 ( .A1(n3357), .A2(reg_file[418]), .B1(n4761), .B2(
        reg_file[386]), .ZN(n5103) );
  AOI22_X1 U6385 ( .A1(n3357), .A2(reg_file[672]), .B1(n4761), .B2(
        reg_file[640]), .ZN(n4984) );
  AOI22_X1 U6386 ( .A1(n3357), .A2(reg_file[160]), .B1(n4761), .B2(
        reg_file[128]), .ZN(n4989) );
  AOI22_X1 U6387 ( .A1(n3357), .A2(reg_file[930]), .B1(n4761), .B2(
        reg_file[898]), .ZN(n5108) );
  AOI22_X1 U6388 ( .A1(n3357), .A2(reg_file[928]), .B1(n4761), .B2(
        reg_file[896]), .ZN(n4994) );
  AOI22_X1 U6389 ( .A1(n3357), .A2(reg_file[161]), .B1(n4761), .B2(
        reg_file[129]), .ZN(n5036) );
  AOI22_X1 U6390 ( .A1(n3357), .A2(reg_file[929]), .B1(n4761), .B2(
        reg_file[897]), .ZN(n5041) );
  AOI22_X1 U6391 ( .A1(n3357), .A2(reg_file[417]), .B1(n4761), .B2(
        reg_file[385]), .ZN(n5046) );
  AOI22_X1 U6392 ( .A1(n3357), .A2(reg_file[673]), .B1(n4761), .B2(
        reg_file[641]), .ZN(n5051) );
  NAND2_X1 U6393 ( .A1(n4965), .A2(n6381), .ZN(n4966) );
  AOI211_X1 U6394 ( .C1(n4824), .C2(rs1_val_gpr_w[1]), .A(n6598), .B(n6893), 
        .ZN(n6599) );
  OAI22_X1 U6395 ( .A1(n4819), .A2(n3825), .B1(n3321), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n98) );
  AOI21_X1 U6396 ( .B1(n6579), .B2(mem_i_inst_i[28]), .A(n6568), .ZN(n6569) );
  OAI22_X1 U6397 ( .A1(n4819), .A2(n3826), .B1(n6548), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n97) );
  OAI22_X1 U6398 ( .A1(n4819), .A2(n3827), .B1(n3379), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n96) );
  OAI22_X1 U6399 ( .A1(n4819), .A2(n3828), .B1(n3306), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n95) );
  OAI22_X1 U6400 ( .A1(n4819), .A2(n3824), .B1(n3324), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n94) );
  AOI21_X1 U6401 ( .B1(n6579), .B2(mem_i_inst_i[11]), .A(n6574), .ZN(n6575) );
  OAI22_X1 U6402 ( .A1(n3287), .A2(n3823), .B1(n3288), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n93) );
  AOI21_X1 U6403 ( .B1(n6579), .B2(mem_i_inst_i[10]), .A(n6578), .ZN(n6580) );
  OAI22_X1 U6404 ( .A1(n3287), .A2(n3771), .B1(n3329), .B2(n3297), .ZN(
        DP_OP_181_135_5161_n92) );
  XNOR2_X1 U6405 ( .A(rs2_val_gpr_w[1]), .B(rs1_val_gpr_w[1]), .ZN(n6430) );
  AOI22_X1 U6406 ( .A1(reg_file[450]), .A2(n4798), .B1(n6383), .B2(
        reg_file[418]), .ZN(n5844) );
  AOI22_X1 U6407 ( .A1(n4798), .A2(reg_file[192]), .B1(n6383), .B2(
        reg_file[160]), .ZN(n4948) );
  AOI22_X1 U6408 ( .A1(n4798), .A2(reg_file[962]), .B1(n6383), .B2(
        reg_file[930]), .ZN(n5849) );
  AOI22_X1 U6409 ( .A1(n4798), .A2(reg_file[194]), .B1(n6383), .B2(
        reg_file[162]), .ZN(n5854) );
  AOI22_X1 U6410 ( .A1(n4798), .A2(reg_file[960]), .B1(n6383), .B2(
        reg_file[928]), .ZN(n4953) );
  AOI22_X1 U6411 ( .A1(n4798), .A2(reg_file[706]), .B1(n6383), .B2(
        reg_file[674]), .ZN(n5859) );
  AOI22_X1 U6412 ( .A1(n4798), .A2(reg_file[704]), .B1(n6383), .B2(
        reg_file[672]), .ZN(n4958) );
  AOI22_X1 U6413 ( .A1(n4798), .A2(reg_file[448]), .B1(n6383), .B2(
        reg_file[416]), .ZN(n4963) );
  AOI22_X1 U6414 ( .A1(n4799), .A2(reg_file[705]), .B1(n6383), .B2(
        reg_file[673]), .ZN(n5820) );
  AOI22_X1 U6415 ( .A1(n4798), .A2(reg_file[961]), .B1(n6383), .B2(
        reg_file[929]), .ZN(n5825) );
  AOI22_X1 U6416 ( .A1(n4798), .A2(reg_file[193]), .B1(n6383), .B2(
        reg_file[161]), .ZN(n5830) );
  AOI22_X1 U6417 ( .A1(n4798), .A2(reg_file[449]), .B1(n6383), .B2(
        reg_file[417]), .ZN(n5835) );
  BUF_X1 U6418 ( .A(n3769), .Z(n4763) );
  BUF_X1 U6419 ( .A(n3769), .Z(n4764) );
  BUF_X1 U6420 ( .A(n3769), .Z(n4765) );
  BUF_X1 U6421 ( .A(n3799), .Z(n4771) );
  BUF_X1 U6422 ( .A(n3799), .Z(n4772) );
  BUF_X1 U6423 ( .A(n3799), .Z(n4773) );
  BUF_X1 U6424 ( .A(n3799), .Z(n4774) );
  BUF_X1 U6425 ( .A(n6383), .Z(n4791) );
  BUF_X1 U6426 ( .A(n6385), .Z(n4803) );
  BUF_X1 U6427 ( .A(n6385), .Z(n4804) );
  XOR2_X1 U6428 ( .A(rs2_val_gpr_w[10]), .B(rs1_val_gpr_w[10]), .Z(n6427) );
  MUX2_X1 U6429 ( .A(n6450), .B(n6854), .S(n6449), .Z(n6453) );
  NAND3_X1 U6430 ( .A1(reset_vector_i[4]), .A2(reset_vector_i[5]), .A3(
        reset_vector_i[6]), .ZN(n6714) );
  INV_X1 U6431 ( .A(reset_vector_i[7]), .ZN(n6713) );
  NOR2_X1 U6432 ( .A1(n6714), .A2(n6713), .ZN(n6712) );
  NAND2_X1 U6433 ( .A1(n6712), .A2(reset_vector_i[8]), .ZN(n6711) );
  INV_X1 U6434 ( .A(reset_vector_i[9]), .ZN(n6710) );
  NOR2_X1 U6435 ( .A1(n6711), .A2(n6710), .ZN(n6709) );
  NAND2_X1 U6436 ( .A1(n6709), .A2(reset_vector_i[10]), .ZN(n6708) );
  INV_X1 U6437 ( .A(reset_vector_i[11]), .ZN(n6707) );
  NOR2_X1 U6438 ( .A1(n6708), .A2(n6707), .ZN(n6706) );
  NAND2_X1 U6439 ( .A1(n6706), .A2(reset_vector_i[12]), .ZN(n6705) );
  INV_X1 U6440 ( .A(reset_vector_i[13]), .ZN(n6704) );
  NOR2_X1 U6441 ( .A1(n6705), .A2(n6704), .ZN(n6703) );
  NAND2_X1 U6442 ( .A1(n6703), .A2(reset_vector_i[14]), .ZN(n6702) );
  INV_X1 U6443 ( .A(reset_vector_i[15]), .ZN(n6701) );
  NOR2_X1 U6444 ( .A1(n6702), .A2(n6701), .ZN(n6700) );
  NAND2_X1 U6445 ( .A1(n6700), .A2(reset_vector_i[16]), .ZN(n6699) );
  INV_X1 U6446 ( .A(reset_vector_i[17]), .ZN(n6698) );
  NOR2_X1 U6447 ( .A1(n6699), .A2(n6698), .ZN(n6697) );
  NAND2_X1 U6448 ( .A1(n6697), .A2(reset_vector_i[18]), .ZN(n6696) );
  INV_X1 U6449 ( .A(reset_vector_i[19]), .ZN(n6695) );
  NOR2_X1 U6450 ( .A1(n6696), .A2(n6695), .ZN(n6694) );
  NAND2_X1 U6451 ( .A1(n6694), .A2(reset_vector_i[20]), .ZN(n6693) );
  INV_X1 U6452 ( .A(reset_vector_i[21]), .ZN(n6692) );
  NOR2_X1 U6453 ( .A1(n6693), .A2(n6692), .ZN(n6691) );
  NAND2_X1 U6454 ( .A1(n6691), .A2(reset_vector_i[22]), .ZN(n6690) );
  INV_X1 U6455 ( .A(reset_vector_i[23]), .ZN(n6689) );
  NOR2_X1 U6456 ( .A1(n6690), .A2(n6689), .ZN(n6688) );
  NAND2_X1 U6457 ( .A1(n6688), .A2(reset_vector_i[24]), .ZN(n6687) );
  XNOR2_X1 U6458 ( .A(n6688), .B(reset_vector_i[24]), .ZN(n6766) );
  AOI21_X1 U6459 ( .B1(n6690), .B2(n6689), .A(n6688), .ZN(n_0_net__23_) );
  XNOR2_X1 U6460 ( .A(n6691), .B(reset_vector_i[22]), .ZN(n6765) );
  XNOR2_X1 U6461 ( .A(n6694), .B(reset_vector_i[20]), .ZN(n6764) );
  AOI21_X1 U6462 ( .B1(n6699), .B2(n6698), .A(n6697), .ZN(n_0_net__17_) );
  XNOR2_X1 U6463 ( .A(n6700), .B(reset_vector_i[16]), .ZN(n6763) );
  AOI21_X1 U6464 ( .B1(n6705), .B2(n6704), .A(n6703), .ZN(n_0_net__13_) );
  XNOR2_X1 U6465 ( .A(n6706), .B(reset_vector_i[12]), .ZN(n6762) );
  XNOR2_X1 U6466 ( .A(n6712), .B(reset_vector_i[8]), .ZN(n6761) );
  INV_X1 U6467 ( .A(reset_vector_i[4]), .ZN(n_0_net__4_) );
  INV_X1 U6468 ( .A(reset_vector_i[5]), .ZN(n6715) );
  NAND3_X1 U6469 ( .A1(n6756), .A2(n6755), .A3(n6754), .ZN(n6758) );
  INV_X1 U6470 ( .A(n6758), .ZN(n6722) );
  NOR3_X1 U6471 ( .A1(n57), .A2(state_q_0_), .A3(n6726), .ZN(n6721) );
  NAND3_X1 U6472 ( .A1(n4910), .A2(n6830), .A3(n6827), .ZN(n6716) );
  NOR3_X1 U6473 ( .A1(mem_i_inst_i[29]), .A2(mem_i_inst_i[28]), .A3(n6716), 
        .ZN(n6729) );
  NAND2_X1 U6474 ( .A1(n6756), .A2(mem_i_inst_i[5]), .ZN(n6717) );
  NAND3_X1 U6475 ( .A1(mem_i_inst_i[4]), .A2(n6686), .A3(n6754), .ZN(n6746) );
  NOR2_X1 U6476 ( .A1(n6717), .A2(n6746), .ZN(n6778) );
  NAND2_X1 U6477 ( .A1(n6729), .A2(n6778), .ZN(n6749) );
  INV_X1 U6478 ( .A(n6721), .ZN(n6720) );
  NOR4_X1 U6479 ( .A1(n57), .A2(state_q_0_), .A3(mem_i_valid_i), .A4(
        muldiv_ready_w), .ZN(n6718) );
  AOI21_X1 U6480 ( .B1(mem_i_rd_o), .B2(mem_i_accept_i), .A(n6718), .ZN(n6719)
         );
  OAI21_X1 U6481 ( .B1(n6743), .B2(n6720), .A(n6719), .ZN(n6725) );
  AOI21_X1 U6482 ( .B1(n6722), .B2(n6721), .A(n6725), .ZN(n6724) );
  NAND2_X1 U6483 ( .A1(state_q_0_), .A2(n3837), .ZN(n6723) );
  AOI221_X1 U6484 ( .B1(mem_d_ack_i), .B2(n6724), .C1(n6723), .C2(n6724), .A(
        rst_i), .ZN(n2917) );
  NOR2_X1 U6485 ( .A1(rst_i), .A2(n6725), .ZN(n2919) );
  NAND2_X1 U6487 ( .A1(n6684), .A2(n6821), .ZN(n6873) );
  NAND4_X1 U6488 ( .A1(mem_i_inst_i[4]), .A2(n6756), .A3(mem_i_inst_i[6]), 
        .A4(mem_i_inst_i[5]), .ZN(n6745) );
  NOR4_X1 U6489 ( .A1(mem_i_inst_i[9]), .A2(mem_i_inst_i[7]), .A3(
        mem_i_inst_i[11]), .A4(mem_i_inst_i[10]), .ZN(n6727) );
  NAND2_X1 U6490 ( .A1(n6727), .A2(n7988), .ZN(n6789) );
  NOR2_X1 U6491 ( .A1(n6745), .A2(n6789), .ZN(n6728) );
  OAI22_X1 U6492 ( .A1(n3331), .A2(rs2_val_gpr_w[27]), .B1(rs1_val_gpr_w[30]), 
        .B2(n3346), .ZN(n6730) );
  OAI22_X1 U6493 ( .A1(n3339), .A2(rs2_val_gpr_w[16]), .B1(rs1_val_gpr_w[22]), 
        .B2(n3343), .ZN(n6731) );
  OAI22_X1 U6494 ( .A1(n3304), .A2(rs2_val_gpr_w[15]), .B1(rs1_val_gpr_w[28]), 
        .B2(n3348), .ZN(n6732) );
  OAI22_X1 U6495 ( .A1(n3289), .A2(rs2_val_gpr_w[11]), .B1(rs1_val_gpr_w[6]), 
        .B2(n3313), .ZN(n6733) );
  OAI22_X1 U6496 ( .A1(n3330), .A2(rs2_val_gpr_w[25]), .B1(rs1_val_gpr_w[7]), 
        .B2(n3292), .ZN(n6734) );
  OAI22_X1 U6497 ( .A1(n3321), .A2(rs2_val_gpr_w[8]), .B1(rs1_val_gpr_w[21]), 
        .B2(n3312), .ZN(n6735) );
  OAI22_X1 U6498 ( .A1(n3308), .A2(rs2_val_gpr_w[9]), .B1(rs1_val_gpr_w[19]), 
        .B2(n3332), .ZN(n6736) );
  OAI22_X1 U6499 ( .A1(n3323), .A2(rs2_val_gpr_w[14]), .B1(rs1_val_gpr_w[13]), 
        .B2(n3291), .ZN(n6737) );
  OAI22_X1 U6500 ( .A1(n3307), .A2(rs2_val_gpr_w[23]), .B1(rs1_val_gpr_w[18]), 
        .B2(n3337), .ZN(n6738) );
  OAI211_X1 U6501 ( .C1(rs2_val_gpr_w[26]), .C2(n3333), .A(n6741), .B(n6740), 
        .ZN(n6739) );
  NOR2_X1 U6502 ( .A1(n6742), .A2(n6743), .ZN(inst_divu_w) );
  AND2_X1 U6503 ( .A1(n6681), .A2(n6750), .ZN(inst_mul_w) );
  NOR2_X1 U6504 ( .A1(n6854), .A2(n6743), .ZN(inst_mulh_w) );
  NOR2_X1 U6505 ( .A1(mem_i_inst_i[14]), .A2(n6684), .ZN(n6783) );
  NAND2_X1 U6506 ( .A1(n6783), .A2(n6685), .ZN(n6855) );
  NOR2_X1 U6507 ( .A1(n6855), .A2(n6743), .ZN(inst_mulhsu_w) );
  AND3_X1 U6508 ( .A1(mem_i_inst_i[12]), .A2(n6783), .A3(n6750), .ZN(
        inst_mulhu_w) );
  NOR3_X1 U6509 ( .A1(mem_i_inst_i[12]), .A2(n6744), .A3(n6743), .ZN(
        inst_rem_w) );
  NOR3_X1 U6510 ( .A1(n6685), .A2(n6744), .A3(n6743), .ZN(inst_remu_w) );
  NOR2_X1 U6511 ( .A1(mem_i_inst_i[5]), .A2(n6758), .ZN(n6844) );
  AOI21_X1 U6512 ( .B1(n6685), .B2(n6684), .A(n6745), .ZN(n6790) );
  INV_X1 U6513 ( .A(mem_i_inst_i[2]), .ZN(n6747) );
  NOR2_X1 U6514 ( .A1(n6747), .A2(n6746), .ZN(n6814) );
  NOR3_X1 U6515 ( .A1(n6679), .A2(n6790), .A3(n6814), .ZN(n6782) );
  NAND4_X1 U6516 ( .A1(n6754), .A2(n6748), .A3(n6756), .A4(mem_i_inst_i[4]), 
        .ZN(n6792) );
  OAI21_X1 U6517 ( .B1(mem_i_inst_i[25]), .B2(n6749), .A(n6792), .ZN(n6776) );
  NOR4_X1 U6518 ( .A1(mem_i_inst_i[5]), .A2(mem_i_inst_i[6]), .A3(n6686), .A4(
        n6873), .ZN(n6751) );
  AOI22_X1 U6519 ( .A1(mem_i_inst_i[2]), .A2(n6751), .B1(n6756), .B2(
        mem_i_inst_i[5]), .ZN(n6752) );
  OAI211_X1 U6520 ( .C1(n6788), .C2(n6753), .A(mem_i_inst_i[0]), .B(
        mem_i_inst_i[1]), .ZN(invalid_inst_r) );
  NAND2_X1 U6521 ( .A1(n6684), .A2(mem_i_inst_i[12]), .ZN(n6872) );
  INV_X1 U6522 ( .A(n6872), .ZN(n6757) );
  NOR2_X1 U6523 ( .A1(n6855), .A2(n6758), .ZN(n6759) );
  AND3_X1 U6524 ( .A1(state_q_0_), .A2(mem_d_ack_i), .A3(n3837), .ZN(n6878) );
  NOR2_X1 U6525 ( .A1(n6878), .A2(muldiv_ready_w), .ZN(n6772) );
  NAND2_X1 U6526 ( .A1(n6877), .A2(n6793), .ZN(n6771) );
  NAND2_X1 U6527 ( .A1(n6683), .A2(n6813), .ZN(n6787) );
  OAI22_X1 U6528 ( .A1(n147), .A2(n6771), .B1(n6787), .B2(n7986), .ZN(n2884)
         );
  OAI22_X1 U6529 ( .A1(n146), .A2(n6771), .B1(n6787), .B2(n7988), .ZN(n2883)
         );
  INV_X1 U6530 ( .A(mem_i_inst_i[9]), .ZN(n7987) );
  OAI22_X1 U6531 ( .A1(n145), .A2(n6771), .B1(n6787), .B2(n7987), .ZN(n2882)
         );
  INV_X1 U6532 ( .A(mem_i_inst_i[10]), .ZN(n7989) );
  OAI22_X1 U6533 ( .A1(n144), .A2(n6771), .B1(n6787), .B2(n7989), .ZN(n2881)
         );
  INV_X1 U6534 ( .A(mem_i_inst_i[11]), .ZN(n7991) );
  OAI22_X1 U6535 ( .A1(n143), .A2(n6771), .B1(n6787), .B2(n7991), .ZN(n2880)
         );
  OAI21_X1 U6536 ( .B1(n6783), .B2(n6685), .A(n6855), .ZN(n6775) );
  AOI221_X1 U6537 ( .B1(mem_i_inst_i[30]), .B2(n6775), .C1(n6774), .C2(n6775), 
        .A(n6682), .ZN(n6777) );
  NAND2_X1 U6538 ( .A1(n6813), .A2(n6776), .ZN(n6784) );
  OAI22_X1 U6539 ( .A1(n157), .A2(n6918), .B1(n6777), .B2(n6784), .ZN(n2879)
         );
  AND3_X1 U6540 ( .A1(mem_i_inst_i[30]), .A2(n6778), .A3(n6685), .ZN(n6779) );
  OAI22_X1 U6541 ( .A1(mem_i_inst_i[12]), .A2(n6821), .B1(n6779), .B2(n6873), 
        .ZN(n6780) );
  OAI22_X1 U6542 ( .A1(n156), .A2(n6918), .B1(n6780), .B2(n6784), .ZN(n2878)
         );
  AOI21_X1 U6543 ( .B1(mem_i_inst_i[12]), .B2(n6680), .A(n6681), .ZN(n6781) );
  OAI222_X1 U6544 ( .A1(n6918), .A2(n155), .B1(n6793), .B2(n6782), .C1(n6784), 
        .C2(n6781), .ZN(n2877) );
  AOI21_X1 U6545 ( .B1(mem_i_inst_i[14]), .B2(n6685), .A(n6783), .ZN(n6785) );
  OAI22_X1 U6546 ( .A1(n154), .A2(n6918), .B1(n6785), .B2(n6784), .ZN(n2876)
         );
  AOI22_X1 U6547 ( .A1(alu_b_q[0]), .A2(n4826), .B1(mem_i_inst_i[20]), .B2(
        n6808), .ZN(n6794) );
  AOI22_X1 U6548 ( .A1(alu_b_q[1]), .A2(n4827), .B1(mem_i_inst_i[21]), .B2(
        n6808), .ZN(n6795) );
  INV_X1 U6549 ( .A(n6808), .ZN(n6811) );
  NAND2_X1 U6550 ( .A1(n6679), .A2(n6813), .ZN(n6879) );
  OAI211_X1 U6551 ( .C1(n3763), .C2(n6918), .A(n6796), .B(n6879), .ZN(n2872)
         );
  AOI22_X1 U6552 ( .A1(alu_b_q[3]), .A2(n4827), .B1(mem_i_inst_i[23]), .B2(
        n6808), .ZN(n6797) );
  AOI22_X1 U6553 ( .A1(alu_b_q[4]), .A2(n4827), .B1(mem_i_inst_i[24]), .B2(
        n6808), .ZN(n6798) );
  AOI22_X1 U6554 ( .A1(alu_b_q[5]), .A2(n4827), .B1(mem_i_inst_i[25]), .B2(
        n6808), .ZN(n6799) );
  AOI22_X1 U6555 ( .A1(csr_data_w[6]), .A2(n6839), .B1(n6840), .B2(
        rs2_val_gpr_w[6]), .ZN(n6801) );
  AOI22_X1 U6556 ( .A1(alu_b_q[6]), .A2(n4827), .B1(mem_i_inst_i[26]), .B2(
        n6808), .ZN(n6800) );
  NAND2_X1 U6557 ( .A1(n6801), .A2(n6800), .ZN(n2868) );
  AOI22_X1 U6558 ( .A1(csr_data_w[7]), .A2(n6839), .B1(n6840), .B2(
        rs2_val_gpr_w[7]), .ZN(n6803) );
  AOI22_X1 U6559 ( .A1(alu_b_q[7]), .A2(n4827), .B1(mem_i_inst_i[27]), .B2(
        n6808), .ZN(n6802) );
  NAND2_X1 U6560 ( .A1(n6803), .A2(n6802), .ZN(n2867) );
  AOI22_X1 U6561 ( .A1(csr_data_w[8]), .A2(n6839), .B1(n6840), .B2(
        rs2_val_gpr_w[8]), .ZN(n6805) );
  AOI22_X1 U6562 ( .A1(alu_b_q[8]), .A2(n4827), .B1(mem_i_inst_i[28]), .B2(
        n6808), .ZN(n6804) );
  NAND2_X1 U6563 ( .A1(n6805), .A2(n6804), .ZN(n2866) );
  AOI22_X1 U6564 ( .A1(csr_data_w[9]), .A2(n6839), .B1(n6840), .B2(
        rs2_val_gpr_w[9]), .ZN(n6807) );
  AOI22_X1 U6565 ( .A1(alu_b_q[9]), .A2(n4827), .B1(mem_i_inst_i[29]), .B2(
        n6808), .ZN(n6806) );
  NAND2_X1 U6566 ( .A1(n6807), .A2(n6806), .ZN(n2865) );
  AOI22_X1 U6567 ( .A1(csr_data_w[10]), .A2(n6839), .B1(n6840), .B2(
        rs2_val_gpr_w[10]), .ZN(n6810) );
  AOI22_X1 U6568 ( .A1(alu_b_q[10]), .A2(n4827), .B1(mem_i_inst_i[30]), .B2(
        n6808), .ZN(n6809) );
  NAND2_X1 U6569 ( .A1(n6810), .A2(n6809), .ZN(n2864) );
  AOI22_X1 U6570 ( .A1(csr_data_w[11]), .A2(n6839), .B1(n6840), .B2(
        rs2_val_gpr_w[11]), .ZN(n6812) );
  OAI211_X1 U6571 ( .C1(n6918), .C2(n3775), .A(n6812), .B(n6841), .ZN(n2863)
         );
  OAI22_X1 U6572 ( .A1(n3350), .A2(n6838), .B1(n6685), .B2(n6880), .ZN(n6815)
         );
  AOI21_X1 U6573 ( .B1(n6839), .B2(csr_data_w[12]), .A(n6815), .ZN(n6816) );
  OAI211_X1 U6574 ( .C1(n6918), .C2(n3806), .A(n6816), .B(n6841), .ZN(n2862)
         );
  OAI22_X1 U6575 ( .A1(n3291), .A2(n6838), .B1(n6684), .B2(n6880), .ZN(n6817)
         );
  AOI21_X1 U6576 ( .B1(n6839), .B2(csr_data_w[13]), .A(n6817), .ZN(n6818) );
  OAI211_X1 U6577 ( .C1(n6918), .C2(n3776), .A(n6818), .B(n6841), .ZN(n2861)
         );
  AOI21_X1 U6578 ( .B1(n4826), .B2(alu_b_q[14]), .A(n6835), .ZN(n6820) );
  AOI22_X1 U6579 ( .A1(csr_data_w[14]), .A2(n6839), .B1(n6840), .B2(
        rs2_val_gpr_w[14]), .ZN(n6819) );
  OAI211_X1 U6580 ( .C1(n6821), .C2(n6880), .A(n6820), .B(n6819), .ZN(n2860)
         );
  AOI21_X1 U6581 ( .B1(n4826), .B2(alu_b_q[25]), .A(n6835), .ZN(n6823) );
  AOI22_X1 U6582 ( .A1(csr_data_w[25]), .A2(n6839), .B1(n6840), .B2(
        rs2_val_gpr_w[25]), .ZN(n6822) );
  OAI211_X1 U6583 ( .C1(n6824), .C2(n6880), .A(n6823), .B(n6822), .ZN(n2849)
         );
  AOI21_X1 U6584 ( .B1(n4826), .B2(alu_b_q[26]), .A(n6835), .ZN(n6826) );
  AOI22_X1 U6585 ( .A1(csr_data_w[26]), .A2(n6839), .B1(n6840), .B2(
        rs2_val_gpr_w[26]), .ZN(n6825) );
  OAI211_X1 U6586 ( .C1(n6827), .C2(n6880), .A(n6826), .B(n6825), .ZN(n2848)
         );
  AOI21_X1 U6587 ( .B1(n4826), .B2(alu_b_q[27]), .A(n6835), .ZN(n6829) );
  AOI22_X1 U6588 ( .A1(csr_data_w[27]), .A2(n6839), .B1(n6840), .B2(
        rs2_val_gpr_w[27]), .ZN(n6828) );
  OAI211_X1 U6589 ( .C1(n6830), .C2(n6880), .A(n6829), .B(n6828), .ZN(n2847)
         );
  AOI21_X1 U6590 ( .B1(n4827), .B2(alu_b_q[28]), .A(n6835), .ZN(n6832) );
  AOI22_X1 U6591 ( .A1(mem_i_inst_i[28]), .A2(n6637), .B1(n6839), .B2(
        csr_data_w[28]), .ZN(n6831) );
  OAI211_X1 U6592 ( .C1(n3348), .C2(n6838), .A(n6832), .B(n6831), .ZN(n2846)
         );
  AOI21_X1 U6593 ( .B1(n4826), .B2(alu_b_q[29]), .A(n6835), .ZN(n6834) );
  AOI22_X1 U6594 ( .A1(csr_data_w[29]), .A2(n6839), .B1(n6840), .B2(
        rs2_val_gpr_w[29]), .ZN(n6833) );
  OAI211_X1 U6595 ( .C1(n6566), .C2(n6880), .A(n6834), .B(n6833), .ZN(n2845)
         );
  AOI21_X1 U6596 ( .B1(n4826), .B2(alu_b_q[30]), .A(n6835), .ZN(n6837) );
  AOI22_X1 U6597 ( .A1(mem_i_inst_i[30]), .A2(n6637), .B1(n6839), .B2(
        csr_data_w[30]), .ZN(n6836) );
  OAI211_X1 U6598 ( .C1(n3346), .C2(n6838), .A(n6837), .B(n6836), .ZN(n2844)
         );
  AOI22_X1 U6599 ( .A1(alu_b_q[31]), .A2(n4827), .B1(n6839), .B2(
        csr_data_w[31]), .ZN(n6843) );
  AOI22_X1 U6600 ( .A1(mem_i_inst_i[31]), .A2(n6637), .B1(n6840), .B2(
        rs2_val_gpr_w[31]), .ZN(n6842) );
  NAND3_X1 U6601 ( .A1(n6843), .A2(n6842), .A3(n6841), .ZN(n2843) );
  NOR2_X1 U6602 ( .A1(mem_d_accept_i), .A2(n3796), .ZN(n6869) );
  AOI22_X1 U6603 ( .A1(n4821), .A2(n6844), .B1(n6869), .B2(mem_d_rd_o), .ZN(
        n1463) );
  NAND2_X1 U6604 ( .A1(n4821), .A2(n7992), .ZN(n6853) );
  NOR2_X1 U6605 ( .A1(n6873), .A2(n6853), .ZN(n6846) );
  NOR2_X1 U6606 ( .A1(n6685), .A2(n6862), .ZN(n6859) );
  AOI22_X1 U6607 ( .A1(n6859), .A2(rs2_val_gpr_w[15]), .B1(n6863), .B2(
        rs2_val_gpr_w[31]), .ZN(n6848) );
  NAND2_X1 U6608 ( .A1(n4822), .A2(mem_d_data_wr_o[31]), .ZN(n6847) );
  OAI211_X1 U6609 ( .C1(n3292), .C2(n6860), .A(n6848), .B(n6847), .ZN(n2842)
         );
  AOI22_X1 U6610 ( .A1(n6859), .A2(rs2_val_gpr_w[14]), .B1(n6863), .B2(
        rs2_val_gpr_w[30]), .ZN(n6850) );
  NAND2_X1 U6611 ( .A1(n4822), .A2(mem_d_data_wr_o[30]), .ZN(n6849) );
  OAI211_X1 U6612 ( .C1(n3313), .C2(n6860), .A(n6850), .B(n6849), .ZN(n2841)
         );
  AOI22_X1 U6613 ( .A1(mem_d_data_wr_o[23]), .A2(n4822), .B1(n6863), .B2(
        rs2_val_gpr_w[23]), .ZN(n6851) );
  OAI21_X1 U6614 ( .B1(n3292), .B2(n6862), .A(n6851), .ZN(n2834) );
  AOI22_X1 U6615 ( .A1(mem_d_data_wr_o[22]), .A2(n4822), .B1(n6863), .B2(
        rs2_val_gpr_w[22]), .ZN(n6852) );
  OAI21_X1 U6616 ( .B1(n3313), .B2(n6862), .A(n6852), .ZN(n2833) );
  AOI22_X1 U6617 ( .A1(mem_d_data_wr_o[15]), .A2(n4822), .B1(rs2_val_gpr_w[15]), .B2(n6677), .ZN(n6856) );
  OAI21_X1 U6618 ( .B1(n3292), .B2(n6865), .A(n6856), .ZN(n2826) );
  AOI22_X1 U6619 ( .A1(mem_d_data_wr_o[14]), .A2(n4822), .B1(rs2_val_gpr_w[14]), .B2(n6677), .ZN(n6857) );
  OAI21_X1 U6620 ( .B1(n3313), .B2(n6865), .A(n6857), .ZN(n2825) );
  AOI22_X1 U6621 ( .A1(mem_d_data_wr_o[7]), .A2(n4822), .B1(rs2_val_gpr_w[7]), 
        .B2(n6868), .ZN(n1387) );
  AOI22_X1 U6622 ( .A1(mem_d_data_wr_o[6]), .A2(n4822), .B1(rs2_val_gpr_w[6]), 
        .B2(n6868), .ZN(n1386) );
  AOI211_X1 U6623 ( .C1(n6869), .C2(mem_d_wr_o[3]), .A(n6863), .B(n6859), .ZN(
        n6861) );
  NAND2_X1 U6624 ( .A1(n6861), .A2(n6860), .ZN(n2818) );
  AOI211_X1 U6625 ( .C1(n6869), .C2(mem_d_wr_o[2]), .A(n6863), .B(n6678), .ZN(
        n6864) );
  INV_X1 U6626 ( .A(n6864), .ZN(n2817) );
  INV_X1 U6627 ( .A(n6869), .ZN(n6867) );
  OAI211_X1 U6628 ( .C1(n6867), .C2(n4708), .A(n6866), .B(n6865), .ZN(n2816)
         );
  AOI21_X1 U6629 ( .B1(n6869), .B2(mem_d_wr_o[0]), .A(n6868), .ZN(n1370) );
  NAND3_X1 U6630 ( .A1(n6870), .A2(n6685), .A3(n6684), .ZN(n6871) );
  OAI21_X1 U6631 ( .B1(n158), .B2(n6875), .A(n6871), .ZN(n2815) );
  OAI22_X1 U6632 ( .A1(n159), .A2(n6875), .B1(n6874), .B2(n6872), .ZN(n2814)
         );
  OAI22_X1 U6633 ( .A1(n162), .A2(n6875), .B1(n6874), .B2(n6873), .ZN(n2811)
         );
  INV_X1 U6634 ( .A(muldiv_ready_w), .ZN(n6876) );
  NAND2_X1 U6635 ( .A1(n6878), .A2(n6877), .ZN(n6883) );
  NOR2_X1 U6636 ( .A1(n158), .A2(n6883), .ZN(n6882) );
  NAND2_X1 U6637 ( .A1(n6882), .A2(n3874), .ZN(n6881) );
  NOR2_X1 U6638 ( .A1(n160), .A2(n6881), .ZN(n6919) );
  AOI22_X1 U6639 ( .A1(n4823), .A2(muldiv_result_w[0]), .B1(n6919), .B2(
        mem_d_data_rd_i[24]), .ZN(n6890) );
  OAI21_X1 U6640 ( .B1(mem_i_inst_i[5]), .B2(n6880), .A(n6879), .ZN(n7008) );
  NOR2_X1 U6641 ( .A1(n3866), .A2(n6881), .ZN(n6920) );
  AOI22_X1 U6642 ( .A1(mem_i_pc_o[0]), .A2(n4825), .B1(n6920), .B2(
        mem_d_data_rd_i[8]), .ZN(n6888) );
  AND2_X1 U6643 ( .A1(n6882), .A2(n161), .ZN(n6921) );
  NAND2_X1 U6644 ( .A1(n6921), .A2(n3866), .ZN(n6885) );
  NOR2_X1 U6645 ( .A1(n160), .A2(n159), .ZN(n6884) );
  NOR2_X1 U6646 ( .A1(n3875), .A2(n6883), .ZN(n6959) );
  NAND2_X1 U6647 ( .A1(n6884), .A2(n6959), .ZN(n6925) );
  NAND2_X1 U6648 ( .A1(n6885), .A2(n6925), .ZN(n6911) );
  NAND2_X1 U6649 ( .A1(n160), .A2(n6921), .ZN(n6886) );
  OAI21_X1 U6650 ( .B1(n160), .B2(n159), .A(n6959), .ZN(n6924) );
  NAND2_X1 U6651 ( .A1(n6886), .A2(n6924), .ZN(n6912) );
  AOI22_X1 U6652 ( .A1(mem_d_data_rd_i[16]), .A2(n6911), .B1(
        mem_d_data_rd_i[0]), .B2(n6912), .ZN(n6887) );
  NAND2_X1 U6653 ( .A1(n6888), .A2(n6887), .ZN(n6889) );
  AOI22_X1 U6654 ( .A1(n6920), .A2(mem_d_data_rd_i[9]), .B1(n4823), .B2(
        muldiv_result_w[1]), .ZN(n6894) );
  AOI22_X1 U6655 ( .A1(mem_d_data_rd_i[25]), .A2(n6919), .B1(
        mem_d_data_rd_i[1]), .B2(n6912), .ZN(n6892) );
  AOI22_X1 U6656 ( .A1(mem_i_pc_o[1]), .A2(n4825), .B1(mem_d_data_rd_i[17]), 
        .B2(n6911), .ZN(n6891) );
  NAND2_X1 U6657 ( .A1(n6892), .A2(n6891), .ZN(n6893) );
  AOI22_X1 U6658 ( .A1(n4823), .A2(muldiv_result_w[2]), .B1(n6919), .B2(
        mem_d_data_rd_i[26]), .ZN(n6898) );
  AOI22_X1 U6659 ( .A1(n6920), .A2(mem_d_data_rd_i[10]), .B1(
        mem_d_data_rd_i[2]), .B2(n6912), .ZN(n6896) );
  AOI22_X1 U6660 ( .A1(mem_i_pc_o[2]), .A2(n4825), .B1(mem_d_data_rd_i[18]), 
        .B2(n6911), .ZN(n6895) );
  NAND2_X1 U6661 ( .A1(n6896), .A2(n6895), .ZN(n6897) );
  AOI22_X1 U6662 ( .A1(n4823), .A2(muldiv_result_w[3]), .B1(n6919), .B2(
        mem_d_data_rd_i[27]), .ZN(n6902) );
  AOI22_X1 U6663 ( .A1(n6920), .A2(mem_d_data_rd_i[11]), .B1(
        mem_d_data_rd_i[19]), .B2(n6911), .ZN(n6900) );
  AOI22_X1 U6664 ( .A1(mem_i_pc_o[3]), .A2(n4825), .B1(mem_d_data_rd_i[3]), 
        .B2(n6912), .ZN(n6899) );
  NAND2_X1 U6665 ( .A1(n6900), .A2(n6899), .ZN(n6901) );
  AOI22_X1 U6666 ( .A1(n6920), .A2(mem_d_data_rd_i[12]), .B1(n4823), .B2(
        muldiv_result_w[4]), .ZN(n6906) );
  AOI22_X1 U6667 ( .A1(mem_d_data_rd_i[28]), .A2(n6919), .B1(
        mem_d_data_rd_i[20]), .B2(n6911), .ZN(n6904) );
  AOI22_X1 U6668 ( .A1(mem_i_pc_o[4]), .A2(n4825), .B1(mem_d_data_rd_i[4]), 
        .B2(n6912), .ZN(n6903) );
  NAND2_X1 U6669 ( .A1(n6904), .A2(n6903), .ZN(n6905) );
  AOI22_X1 U6670 ( .A1(n6920), .A2(mem_d_data_rd_i[13]), .B1(n4823), .B2(
        muldiv_result_w[5]), .ZN(n6910) );
  AOI22_X1 U6671 ( .A1(mem_d_data_rd_i[29]), .A2(n6919), .B1(
        mem_d_data_rd_i[21]), .B2(n6911), .ZN(n6908) );
  AOI22_X1 U6672 ( .A1(mem_i_pc_o[5]), .A2(n4825), .B1(mem_d_data_rd_i[5]), 
        .B2(n6912), .ZN(n6907) );
  NAND2_X1 U6673 ( .A1(n6908), .A2(n6907), .ZN(n6909) );
  AOI22_X1 U6674 ( .A1(n6920), .A2(mem_d_data_rd_i[14]), .B1(n4823), .B2(
        muldiv_result_w[6]), .ZN(n6917) );
  AOI22_X1 U6675 ( .A1(mem_d_data_rd_i[30]), .A2(n6919), .B1(
        mem_d_data_rd_i[22]), .B2(n6911), .ZN(n6914) );
  AOI22_X1 U6676 ( .A1(mem_i_pc_o[6]), .A2(n4825), .B1(mem_d_data_rd_i[6]), 
        .B2(n6912), .ZN(n6913) );
  NAND2_X1 U6677 ( .A1(n6914), .A2(n6913), .ZN(n6915) );
  AOI21_X1 U6678 ( .B1(n4824), .B2(rs1_val_gpr_w[6]), .A(n6915), .ZN(n6916) );
  OAI211_X1 U6679 ( .C1(n3773), .C2(n6918), .A(n6917), .B(n6916), .ZN(n2804)
         );
  AOI22_X1 U6680 ( .A1(n6920), .A2(mem_d_data_rd_i[15]), .B1(n6919), .B2(
        mem_d_data_rd_i[31]), .ZN(n6923) );
  OAI221_X1 U6681 ( .B1(n160), .B2(mem_d_data_rd_i[23]), .C1(n3866), .C2(
        mem_d_data_rd_i[7]), .A(n6921), .ZN(n6922) );
  NAND2_X1 U6682 ( .A1(n6923), .A2(n6922), .ZN(n6958) );
  INV_X1 U6683 ( .A(n6958), .ZN(n6929) );
  AOI22_X1 U6684 ( .A1(alu_a_q[7]), .A2(n4827), .B1(n4823), .B2(
        muldiv_result_w[7]), .ZN(n6928) );
  AOI22_X1 U6685 ( .A1(n6952), .A2(mem_d_data_rd_i[7]), .B1(n6951), .B2(
        mem_d_data_rd_i[23]), .ZN(n6927) );
  AOI22_X1 U6686 ( .A1(mem_i_pc_o[7]), .A2(n4825), .B1(n4824), .B2(n3523), 
        .ZN(n6926) );
  NAND4_X1 U6687 ( .A1(n6929), .A2(n6928), .A3(n6927), .A4(n6926), .ZN(n2803)
         );
  AOI22_X1 U6688 ( .A1(n6951), .A2(mem_d_data_rd_i[24]), .B1(n4823), .B2(
        muldiv_result_w[8]), .ZN(n6932) );
  AOI22_X1 U6689 ( .A1(alu_a_q[8]), .A2(n4827), .B1(mem_d_data_rd_i[8]), .B2(
        n6952), .ZN(n6931) );
  AOI22_X1 U6690 ( .A1(mem_i_pc_o[8]), .A2(n4825), .B1(n4824), .B2(
        rs1_val_gpr_w[8]), .ZN(n6930) );
  NAND2_X1 U6691 ( .A1(n3867), .A2(n6958), .ZN(n6953) );
  NAND4_X1 U6692 ( .A1(n6932), .A2(n6931), .A3(n6930), .A4(n6953), .ZN(n2802)
         );
  AOI22_X1 U6693 ( .A1(alu_a_q[9]), .A2(n4827), .B1(n6952), .B2(
        mem_d_data_rd_i[9]), .ZN(n6935) );
  AOI22_X1 U6694 ( .A1(n6951), .A2(mem_d_data_rd_i[25]), .B1(n4823), .B2(
        muldiv_result_w[9]), .ZN(n6934) );
  AOI22_X1 U6695 ( .A1(mem_i_pc_o[9]), .A2(n4825), .B1(n7007), .B2(
        rs1_val_gpr_w[9]), .ZN(n6933) );
  NAND4_X1 U6696 ( .A1(n6935), .A2(n6934), .A3(n6933), .A4(n6953), .ZN(n2801)
         );
  AOI22_X1 U6697 ( .A1(n6951), .A2(mem_d_data_rd_i[26]), .B1(n4823), .B2(
        muldiv_result_w[10]), .ZN(n6938) );
  AOI22_X1 U6698 ( .A1(alu_a_q[10]), .A2(n4827), .B1(n6952), .B2(
        mem_d_data_rd_i[10]), .ZN(n6937) );
  AOI22_X1 U6699 ( .A1(mem_i_pc_o[10]), .A2(n4825), .B1(n4824), .B2(
        rs1_val_gpr_w[10]), .ZN(n6936) );
  NAND4_X1 U6700 ( .A1(n6938), .A2(n6937), .A3(n6936), .A4(n6953), .ZN(n2800)
         );
  AOI22_X1 U6701 ( .A1(alu_a_q[11]), .A2(n4827), .B1(n6952), .B2(
        mem_d_data_rd_i[11]), .ZN(n6941) );
  AOI22_X1 U6702 ( .A1(n6951), .A2(mem_d_data_rd_i[27]), .B1(n4823), .B2(
        muldiv_result_w[11]), .ZN(n6940) );
  AOI22_X1 U6703 ( .A1(mem_i_pc_o[11]), .A2(n7008), .B1(n4824), .B2(
        rs1_val_gpr_w[11]), .ZN(n6939) );
  NAND4_X1 U6704 ( .A1(n6941), .A2(n6940), .A3(n6939), .A4(n6953), .ZN(n2799)
         );
  AOI22_X1 U6705 ( .A1(alu_a_q[12]), .A2(n4827), .B1(n6952), .B2(
        mem_d_data_rd_i[12]), .ZN(n6944) );
  AOI22_X1 U6706 ( .A1(n6951), .A2(mem_d_data_rd_i[28]), .B1(n4823), .B2(
        muldiv_result_w[12]), .ZN(n6943) );
  AOI22_X1 U6707 ( .A1(mem_i_pc_o[12]), .A2(n7008), .B1(n4824), .B2(
        rs1_val_gpr_w[12]), .ZN(n6942) );
  NAND4_X1 U6708 ( .A1(n6944), .A2(n6943), .A3(n6942), .A4(n6953), .ZN(n2798)
         );
  AOI22_X1 U6709 ( .A1(n6951), .A2(mem_d_data_rd_i[29]), .B1(n7006), .B2(
        muldiv_result_w[13]), .ZN(n6947) );
  AOI22_X1 U6710 ( .A1(alu_a_q[13]), .A2(n4827), .B1(n6952), .B2(
        mem_d_data_rd_i[13]), .ZN(n6946) );
  AOI22_X1 U6711 ( .A1(mem_i_pc_o[13]), .A2(n7008), .B1(n4824), .B2(
        rs1_val_gpr_w[13]), .ZN(n6945) );
  NAND4_X1 U6712 ( .A1(n6947), .A2(n6946), .A3(n6945), .A4(n6953), .ZN(n2797)
         );
  AOI22_X1 U6713 ( .A1(n6951), .A2(mem_d_data_rd_i[30]), .B1(n4823), .B2(
        muldiv_result_w[14]), .ZN(n6950) );
  AOI22_X1 U6714 ( .A1(alu_a_q[14]), .A2(n4827), .B1(n6952), .B2(
        mem_d_data_rd_i[14]), .ZN(n6949) );
  AOI22_X1 U6715 ( .A1(mem_i_pc_o[14]), .A2(n7008), .B1(n4824), .B2(
        rs1_val_gpr_w[14]), .ZN(n6948) );
  NAND4_X1 U6716 ( .A1(n6950), .A2(n6949), .A3(n6948), .A4(n6953), .ZN(n2796)
         );
  AOI22_X1 U6717 ( .A1(n6952), .A2(mem_d_data_rd_i[15]), .B1(n6951), .B2(
        mem_d_data_rd_i[31]), .ZN(n6956) );
  AOI22_X1 U6718 ( .A1(alu_a_q[15]), .A2(n4827), .B1(n7006), .B2(
        muldiv_result_w[15]), .ZN(n6955) );
  AOI22_X1 U6719 ( .A1(mem_i_pc_o[15]), .A2(n7008), .B1(n4824), .B2(
        rs1_val_gpr_w[15]), .ZN(n6954) );
  NAND4_X1 U6720 ( .A1(n6956), .A2(n6955), .A3(n6954), .A4(n6953), .ZN(n2795)
         );
  NOR2_X1 U6721 ( .A1(n6956), .A2(n159), .ZN(n6957) );
  AOI22_X1 U6722 ( .A1(alu_a_q[16]), .A2(n4826), .B1(mem_d_data_rd_i[16]), 
        .B2(n7005), .ZN(n6962) );
  AOI22_X1 U6723 ( .A1(mem_i_pc_o[16]), .A2(n7008), .B1(n4824), .B2(
        rs1_val_gpr_w[16]), .ZN(n6961) );
  NAND2_X1 U6724 ( .A1(n4823), .A2(muldiv_result_w[16]), .ZN(n6960) );
  NAND4_X1 U6725 ( .A1(n7012), .A2(n6962), .A3(n6961), .A4(n6960), .ZN(n2794)
         );
  AOI22_X1 U6726 ( .A1(n7006), .A2(muldiv_result_w[17]), .B1(
        mem_d_data_rd_i[17]), .B2(n7005), .ZN(n6965) );
  AOI22_X1 U6727 ( .A1(mem_i_pc_o[17]), .A2(n7008), .B1(n4824), .B2(
        rs1_val_gpr_w[17]), .ZN(n6964) );
  NAND2_X1 U6728 ( .A1(alu_a_q[17]), .A2(n4826), .ZN(n6963) );
  NAND4_X1 U6729 ( .A1(n7012), .A2(n6965), .A3(n6964), .A4(n6963), .ZN(n2793)
         );
  AOI22_X1 U6730 ( .A1(n4823), .A2(muldiv_result_w[18]), .B1(
        mem_d_data_rd_i[18]), .B2(n7005), .ZN(n6968) );
  AOI22_X1 U6731 ( .A1(mem_i_pc_o[18]), .A2(n7008), .B1(n4824), .B2(
        rs1_val_gpr_w[18]), .ZN(n6967) );
  NAND2_X1 U6732 ( .A1(alu_a_q[18]), .A2(n4827), .ZN(n6966) );
  NAND4_X1 U6733 ( .A1(n7012), .A2(n6968), .A3(n6967), .A4(n6966), .ZN(n2792)
         );
  AOI22_X1 U6734 ( .A1(alu_a_q[19]), .A2(n4827), .B1(mem_d_data_rd_i[19]), 
        .B2(n7005), .ZN(n6971) );
  AOI22_X1 U6735 ( .A1(mem_i_pc_o[19]), .A2(n7008), .B1(n4824), .B2(
        rs1_val_gpr_w[19]), .ZN(n6970) );
  NAND2_X1 U6736 ( .A1(n4823), .A2(muldiv_result_w[19]), .ZN(n6969) );
  NAND4_X1 U6737 ( .A1(n7012), .A2(n6971), .A3(n6970), .A4(n6969), .ZN(n2791)
         );
  AOI22_X1 U6738 ( .A1(n7006), .A2(muldiv_result_w[20]), .B1(
        mem_d_data_rd_i[20]), .B2(n7005), .ZN(n6974) );
  AOI22_X1 U6739 ( .A1(mem_i_pc_o[20]), .A2(n7008), .B1(n4824), .B2(
        rs1_val_gpr_w[20]), .ZN(n6973) );
  NAND2_X1 U6740 ( .A1(alu_a_q[20]), .A2(n4827), .ZN(n6972) );
  NAND4_X1 U6741 ( .A1(n7012), .A2(n6974), .A3(n6973), .A4(n6972), .ZN(n2790)
         );
  AOI22_X1 U6742 ( .A1(alu_a_q[21]), .A2(n4826), .B1(mem_d_data_rd_i[21]), 
        .B2(n7005), .ZN(n6977) );
  AOI22_X1 U6743 ( .A1(mem_i_pc_o[21]), .A2(n7008), .B1(n4824), .B2(
        rs1_val_gpr_w[21]), .ZN(n6976) );
  NAND2_X1 U6744 ( .A1(n4823), .A2(muldiv_result_w[21]), .ZN(n6975) );
  NAND4_X1 U6745 ( .A1(n7012), .A2(n6977), .A3(n6976), .A4(n6975), .ZN(n2789)
         );
  AOI22_X1 U6746 ( .A1(n7006), .A2(muldiv_result_w[22]), .B1(
        mem_d_data_rd_i[22]), .B2(n7005), .ZN(n6980) );
  AOI22_X1 U6747 ( .A1(mem_i_pc_o[22]), .A2(n4825), .B1(n4824), .B2(
        rs1_val_gpr_w[22]), .ZN(n6979) );
  NAND2_X1 U6748 ( .A1(alu_a_q[22]), .A2(n4826), .ZN(n6978) );
  NAND4_X1 U6749 ( .A1(n7012), .A2(n6980), .A3(n6979), .A4(n6978), .ZN(n2788)
         );
  AOI22_X1 U6750 ( .A1(n7006), .A2(muldiv_result_w[23]), .B1(
        mem_d_data_rd_i[23]), .B2(n7005), .ZN(n6983) );
  AOI22_X1 U6751 ( .A1(mem_i_pc_o[23]), .A2(n4825), .B1(n4824), .B2(
        rs1_val_gpr_w[23]), .ZN(n6982) );
  NAND2_X1 U6752 ( .A1(alu_a_q[23]), .A2(n4827), .ZN(n6981) );
  NAND4_X1 U6753 ( .A1(n7012), .A2(n6983), .A3(n6982), .A4(n6981), .ZN(n2787)
         );
  AOI22_X1 U6754 ( .A1(alu_a_q[24]), .A2(n4826), .B1(mem_d_data_rd_i[24]), 
        .B2(n7005), .ZN(n6986) );
  AOI22_X1 U6755 ( .A1(mem_i_pc_o[24]), .A2(n4825), .B1(n4824), .B2(
        rs1_val_gpr_w[24]), .ZN(n6985) );
  NAND2_X1 U6756 ( .A1(n4823), .A2(muldiv_result_w[24]), .ZN(n6984) );
  NAND4_X1 U6757 ( .A1(n7012), .A2(n6986), .A3(n6985), .A4(n6984), .ZN(n2786)
         );
  AOI22_X1 U6758 ( .A1(alu_a_q[25]), .A2(n4826), .B1(mem_d_data_rd_i[25]), 
        .B2(n7005), .ZN(n6989) );
  AOI22_X1 U6759 ( .A1(mem_i_pc_o[25]), .A2(n4825), .B1(n4824), .B2(
        rs1_val_gpr_w[25]), .ZN(n6988) );
  NAND2_X1 U6760 ( .A1(n4823), .A2(muldiv_result_w[25]), .ZN(n6987) );
  NAND4_X1 U6761 ( .A1(n7012), .A2(n6989), .A3(n6988), .A4(n6987), .ZN(n2785)
         );
  AOI22_X1 U6762 ( .A1(alu_a_q[26]), .A2(n4826), .B1(mem_d_data_rd_i[26]), 
        .B2(n7005), .ZN(n6992) );
  NAND2_X1 U6763 ( .A1(n4823), .A2(muldiv_result_w[26]), .ZN(n6990) );
  NAND4_X1 U6764 ( .A1(n7012), .A2(n6992), .A3(n6991), .A4(n6990), .ZN(n2784)
         );
  AOI22_X1 U6765 ( .A1(alu_a_q[27]), .A2(n4826), .B1(mem_d_data_rd_i[27]), 
        .B2(n7005), .ZN(n6995) );
  NAND2_X1 U6766 ( .A1(n4823), .A2(muldiv_result_w[27]), .ZN(n6993) );
  NAND4_X1 U6767 ( .A1(n7012), .A2(n6995), .A3(n6994), .A4(n6993), .ZN(n2783)
         );
  AOI22_X1 U6768 ( .A1(alu_a_q[28]), .A2(n4826), .B1(mem_d_data_rd_i[28]), 
        .B2(n7005), .ZN(n6998) );
  NAND2_X1 U6769 ( .A1(n4823), .A2(muldiv_result_w[28]), .ZN(n6996) );
  NAND4_X1 U6770 ( .A1(n7012), .A2(n6998), .A3(n6997), .A4(n6996), .ZN(n2782)
         );
  AOI22_X1 U6771 ( .A1(alu_a_q[29]), .A2(n4826), .B1(mem_d_data_rd_i[29]), 
        .B2(n7005), .ZN(n7001) );
  NAND2_X1 U6772 ( .A1(n4823), .A2(muldiv_result_w[29]), .ZN(n6999) );
  NAND4_X1 U6773 ( .A1(n7012), .A2(n7001), .A3(n7000), .A4(n6999), .ZN(n2781)
         );
  AOI22_X1 U6774 ( .A1(alu_a_q[30]), .A2(n4826), .B1(mem_d_data_rd_i[30]), 
        .B2(n7005), .ZN(n7004) );
  NAND2_X1 U6775 ( .A1(n4823), .A2(muldiv_result_w[30]), .ZN(n7002) );
  NAND4_X1 U6776 ( .A1(n7012), .A2(n7004), .A3(n7003), .A4(n7002), .ZN(n2780)
         );
  AOI22_X1 U6777 ( .A1(n7006), .A2(muldiv_result_w[31]), .B1(
        mem_d_data_rd_i[31]), .B2(n7005), .ZN(n7011) );
  NAND2_X1 U6778 ( .A1(alu_a_q[31]), .A2(n4826), .ZN(n7009) );
  NAND4_X1 U6779 ( .A1(n7012), .A2(n7011), .A3(n7010), .A4(n7009), .ZN(n2779)
         );
  NOR2_X1 U6780 ( .A1(n3833), .A2(n7082), .ZN(n7838) );
  AOI21_X1 U6781 ( .B1(n7125), .B2(alu_a_q[31]), .A(n7838), .ZN(n7013) );
  NAND2_X1 U6782 ( .A1(n3830), .A2(alu_a_q[31]), .ZN(n7429) );
  INV_X1 U6783 ( .A(n7429), .ZN(n7857) );
  NAND2_X1 U6784 ( .A1(alu_b_q[1]), .A2(n7857), .ZN(n7057) );
  OAI211_X1 U6785 ( .C1(n7774), .C2(n3797), .A(n7013), .B(n7057), .ZN(n7316)
         );
  NOR2_X1 U6786 ( .A1(n3795), .A2(n7082), .ZN(n7599) );
  NOR2_X1 U6787 ( .A1(n3789), .A2(n7122), .ZN(n7703) );
  NOR2_X1 U6788 ( .A1(n3792), .A2(n7883), .ZN(n7649) );
  NOR2_X1 U6789 ( .A1(n3766), .A2(n7774), .ZN(n7550) );
  NOR4_X1 U6790 ( .A1(n7599), .A2(n7703), .A3(n7649), .A4(n7550), .ZN(n7307)
         );
  NOR2_X1 U6791 ( .A1(n7307), .A2(n7282), .ZN(n7015) );
  NOR2_X1 U6792 ( .A1(n3832), .A2(n7082), .ZN(n7704) );
  NOR2_X1 U6793 ( .A1(n3790), .A2(n7122), .ZN(n7836) );
  NOR2_X1 U6794 ( .A1(n3829), .A2(n7774), .ZN(n7652) );
  NOR2_X1 U6795 ( .A1(n3784), .A2(n7883), .ZN(n7777) );
  NOR4_X1 U6796 ( .A1(n7704), .A2(n7836), .A3(n7652), .A4(n7777), .ZN(n7322)
         );
  NOR2_X1 U6797 ( .A1(n3791), .A2(n7122), .ZN(n7600) );
  NOR2_X1 U6798 ( .A1(n3786), .A2(n7082), .ZN(n7502) );
  NOR2_X1 U6799 ( .A1(n3787), .A2(n7883), .ZN(n7548) );
  NOR2_X1 U6800 ( .A1(n3794), .A2(n7774), .ZN(n7448) );
  NOR4_X1 U6801 ( .A1(n7600), .A2(n7502), .A3(n7548), .A4(n7448), .ZN(n7306)
         );
  OAI22_X1 U6802 ( .A1(n7322), .A2(n7313), .B1(n7306), .B2(n7427), .ZN(n7014)
         );
  AOI211_X1 U6803 ( .C1(n7418), .C2(n7316), .A(n7015), .B(n7014), .ZN(n7464)
         );
  INV_X1 U6804 ( .A(n7418), .ZN(n7379) );
  NOR2_X1 U6805 ( .A1(n7379), .A2(alu_b_q[4]), .ZN(n7077) );
  NOR2_X1 U6806 ( .A1(n3793), .A2(n7122), .ZN(n7501) );
  NOR2_X1 U6807 ( .A1(n3785), .A2(n7883), .ZN(n7449) );
  NOR2_X1 U6808 ( .A1(n7501), .A2(n7449), .ZN(n7016) );
  NAND2_X1 U6809 ( .A1(alu_a_q[14]), .A2(n7101), .ZN(n7376) );
  NAND2_X1 U6810 ( .A1(alu_a_q[13]), .A2(n7743), .ZN(n7310) );
  NAND3_X1 U6811 ( .A1(n7016), .A2(n7376), .A3(n7310), .ZN(n7319) );
  NOR2_X1 U6812 ( .A1(n7427), .A2(alu_b_q[4]), .ZN(n7748) );
  NAND2_X1 U6813 ( .A1(alu_a_q[2]), .A2(n7101), .ZN(n7070) );
  NAND2_X1 U6814 ( .A1(alu_a_q[4]), .A2(n7146), .ZN(n7172) );
  NAND2_X1 U6815 ( .A1(alu_a_q[1]), .A2(n7743), .ZN(n7018) );
  NAND2_X1 U6816 ( .A1(alu_a_q[3]), .A2(n7125), .ZN(n7017) );
  NAND4_X1 U6817 ( .A1(n7070), .A2(n7172), .A3(n7018), .A4(n7017), .ZN(n7019)
         );
  AOI22_X1 U6818 ( .A1(n7077), .A2(n7319), .B1(n7748), .B2(n7019), .ZN(n7022)
         );
  NOR2_X1 U6819 ( .A1(n7313), .A2(alu_b_q[4]), .ZN(n7749) );
  NAND2_X1 U6820 ( .A1(alu_a_q[12]), .A2(n7146), .ZN(n7374) );
  NAND2_X1 U6821 ( .A1(alu_a_q[10]), .A2(n7101), .ZN(n7265) );
  NAND2_X1 U6822 ( .A1(alu_a_q[9]), .A2(n7743), .ZN(n7215) );
  NAND2_X1 U6823 ( .A1(alu_a_q[11]), .A2(n7125), .ZN(n7311) );
  NAND4_X1 U6824 ( .A1(n7374), .A2(n7265), .A3(n7215), .A4(n7311), .ZN(n7220)
         );
  NOR2_X1 U6825 ( .A1(n7282), .A2(alu_b_q[4]), .ZN(n7740) );
  NAND2_X1 U6826 ( .A1(alu_a_q[8]), .A2(n7146), .ZN(n7266) );
  NAND2_X1 U6827 ( .A1(alu_a_q[6]), .A2(n7101), .ZN(n7170) );
  NAND2_X1 U6828 ( .A1(alu_a_q[5]), .A2(n7743), .ZN(n7020) );
  NAND2_X1 U6829 ( .A1(alu_a_q[7]), .A2(n7125), .ZN(n7216) );
  NAND4_X1 U6830 ( .A1(n7266), .A2(n7170), .A3(n7020), .A4(n7216), .ZN(n7127)
         );
  AOI22_X1 U6831 ( .A1(n7749), .A2(n7220), .B1(n7740), .B2(n7127), .ZN(n7021)
         );
  OAI211_X1 U6832 ( .C1(n7464), .C2(n3809), .A(n7022), .B(n7021), .ZN(n7033)
         );
  INV_X1 U6833 ( .A(n7068), .ZN(n7876) );
  AOI22_X1 U6834 ( .A1(n3352), .A2(n7876), .B1(n3353), .B2(n7870), .ZN(n7030)
         );
  NAND3_X1 U6835 ( .A1(n3765), .A2(n3788), .A3(n154), .ZN(n7660) );
  NAND2_X1 U6836 ( .A1(n7788), .A2(n7734), .ZN(n7342) );
  NOR2_X1 U6837 ( .A1(n3779), .A2(n7342), .ZN(n7024) );
  OAI22_X1 U6838 ( .A1(n7876), .A2(n3764), .B1(n7870), .B2(n3842), .ZN(n7026)
         );
  NOR3_X1 U6839 ( .A1(n7624), .A2(alu_a_q[1]), .A3(n7026), .ZN(n7023) );
  AOI211_X1 U6840 ( .C1(n7030), .C2(n7024), .A(n7023), .B(n3807), .ZN(n7032)
         );
  NAND2_X1 U6841 ( .A1(n3807), .A2(n3779), .ZN(n7029) );
  NAND2_X1 U6842 ( .A1(n3830), .A2(n155), .ZN(n7025) );
  OAI22_X1 U6843 ( .A1(n3779), .A2(n7774), .B1(n3808), .B2(n7082), .ZN(n7446)
         );
  AOI22_X1 U6844 ( .A1(alu_a_q[1]), .A2(n7802), .B1(n7866), .B2(n7446), .ZN(
        n7028) );
  OAI21_X1 U6845 ( .B1(n7835), .B2(n7026), .A(n7048), .ZN(n7027) );
  OAI211_X1 U6846 ( .C1(n7030), .C2(n7029), .A(n7028), .B(n7027), .ZN(n7031)
         );
  NOR2_X1 U6847 ( .A1(n3807), .A2(n3779), .ZN(n7049) );
  INV_X1 U6848 ( .A(n7073), .ZN(n7050) );
  AOI22_X1 U6849 ( .A1(n3352), .A2(n7071), .B1(n3353), .B2(n7050), .ZN(n7053)
         );
  OAI221_X1 U6850 ( .B1(n3803), .B2(n7053), .C1(n3803), .C2(n7788), .A(n7734), 
        .ZN(n7067) );
  NAND2_X1 U6851 ( .A1(n3763), .A2(n3803), .ZN(n7054) );
  OAI22_X1 U6852 ( .A1(n7050), .A2(n3842), .B1(n3764), .B2(n7071), .ZN(n7051)
         );
  OAI22_X1 U6853 ( .A1(n7835), .A2(n7051), .B1(n3803), .B2(n3763), .ZN(n7055)
         );
  NAND2_X1 U6854 ( .A1(alu_a_q[1]), .A2(n7101), .ZN(n7881) );
  NAND2_X1 U6855 ( .A1(alu_a_q[2]), .A2(n7743), .ZN(n7061) );
  OAI211_X1 U6856 ( .C1(n7883), .C2(n3808), .A(n7881), .B(n7061), .ZN(n7478)
         );
  AOI22_X1 U6857 ( .A1(alu_a_q[2]), .A2(n7802), .B1(n7866), .B2(n7478), .ZN(
        n7052) );
  OAI221_X1 U6858 ( .B1(n7074), .B2(n7055), .C1(n7054), .C2(n7053), .A(n7052), 
        .ZN(n7066) );
  NAND2_X1 U6859 ( .A1(alu_a_q[22]), .A2(n7743), .ZN(n7568) );
  NAND2_X1 U6860 ( .A1(alu_a_q[24]), .A2(n7125), .ZN(n7673) );
  NAND2_X1 U6861 ( .A1(alu_a_q[25]), .A2(n7146), .ZN(n7744) );
  NAND2_X1 U6862 ( .A1(alu_a_q[23]), .A2(n7101), .ZN(n7616) );
  NAND4_X1 U6863 ( .A1(n7568), .A2(n7673), .A3(n7744), .A4(n7616), .ZN(n7355)
         );
  NAND2_X1 U6864 ( .A1(alu_a_q[28]), .A2(n7125), .ZN(n7803) );
  NAND2_X1 U6865 ( .A1(alu_a_q[26]), .A2(n7743), .ZN(n7672) );
  NAND2_X1 U6866 ( .A1(alu_a_q[27]), .A2(n7101), .ZN(n7745) );
  NAND3_X1 U6867 ( .A1(n7803), .A2(n7672), .A3(n7745), .ZN(n7056) );
  AOI21_X1 U6868 ( .B1(alu_a_q[29]), .B2(n7146), .A(n7056), .ZN(n7352) );
  NAND2_X1 U6869 ( .A1(alu_a_q[20]), .A2(n7125), .ZN(n7569) );
  NAND2_X1 U6870 ( .A1(alu_a_q[18]), .A2(n7743), .ZN(n7474) );
  NAND2_X1 U6871 ( .A1(alu_a_q[19]), .A2(n7101), .ZN(n7523) );
  NAND2_X1 U6872 ( .A1(alu_a_q[21]), .A2(n7146), .ZN(n7615) );
  NAND4_X1 U6873 ( .A1(n7569), .A2(n7474), .A3(n7523), .A4(n7615), .ZN(n7357)
         );
  NAND2_X1 U6874 ( .A1(alu_a_q[30]), .A2(n7743), .ZN(n7806) );
  OAI211_X1 U6875 ( .C1(n7082), .C2(n3831), .A(n7806), .B(n7057), .ZN(n7341)
         );
  AOI22_X1 U6876 ( .A1(n7414), .A2(n7357), .B1(n7418), .B2(n7341), .ZN(n7058)
         );
  OAI21_X1 U6877 ( .B1(n7352), .B2(n7313), .A(n7058), .ZN(n7059) );
  AOI21_X1 U6878 ( .B1(n7424), .B2(n7355), .A(n7059), .ZN(n7486) );
  NAND2_X1 U6879 ( .A1(n7699), .A2(n7414), .ZN(n7389) );
  NAND2_X1 U6880 ( .A1(alu_a_q[4]), .A2(n7125), .ZN(n7147) );
  NAND2_X1 U6881 ( .A1(alu_a_q[3]), .A2(n7101), .ZN(n7060) );
  NAND2_X1 U6882 ( .A1(alu_a_q[5]), .A2(n7146), .ZN(n7190) );
  NAND4_X1 U6883 ( .A1(n7147), .A2(n7061), .A3(n7060), .A4(n7190), .ZN(n7062)
         );
  NAND2_X1 U6884 ( .A1(n7699), .A2(n7418), .ZN(n7383) );
  INV_X1 U6885 ( .A(n7383), .ZN(n7354) );
  NAND2_X1 U6886 ( .A1(alu_a_q[16]), .A2(n7125), .ZN(n7475) );
  NAND2_X1 U6887 ( .A1(alu_a_q[14]), .A2(n7743), .ZN(n7346) );
  NAND2_X1 U6888 ( .A1(alu_a_q[17]), .A2(n7146), .ZN(n7522) );
  NAND2_X1 U6889 ( .A1(alu_a_q[15]), .A2(n7101), .ZN(n7421) );
  NAND4_X1 U6890 ( .A1(n7475), .A2(n7346), .A3(n7522), .A4(n7421), .ZN(n7358)
         );
  AOI22_X1 U6891 ( .A1(n7885), .A2(n7062), .B1(n7354), .B2(n7358), .ZN(n7064)
         );
  NAND2_X1 U6892 ( .A1(n7699), .A2(n7424), .ZN(n7385) );
  NAND2_X1 U6893 ( .A1(alu_a_q[6]), .A2(n7743), .ZN(n7148) );
  NAND2_X1 U6894 ( .A1(alu_a_q[8]), .A2(n7125), .ZN(n7229) );
  NAND2_X1 U6895 ( .A1(alu_a_q[9]), .A2(n7146), .ZN(n7276) );
  NAND2_X1 U6896 ( .A1(alu_a_q[7]), .A2(n7101), .ZN(n7189) );
  NAND4_X1 U6897 ( .A1(n7148), .A2(n7229), .A3(n7276), .A4(n7189), .ZN(n7150)
         );
  NOR2_X1 U6898 ( .A1(n7831), .A2(n7313), .ZN(n7356) );
  NAND2_X1 U6899 ( .A1(alu_a_q[10]), .A2(n7743), .ZN(n7228) );
  NAND2_X1 U6900 ( .A1(alu_a_q[12]), .A2(n7125), .ZN(n7345) );
  NAND2_X1 U6901 ( .A1(alu_a_q[13]), .A2(n7146), .ZN(n7420) );
  NAND2_X1 U6902 ( .A1(alu_a_q[11]), .A2(n7101), .ZN(n7277) );
  NAND4_X1 U6903 ( .A1(n7228), .A2(n7345), .A3(n7420), .A4(n7277), .ZN(n7234)
         );
  AOI22_X1 U6904 ( .A1(n7874), .A2(n7150), .B1(n7356), .B2(n7234), .ZN(n7063)
         );
  OAI211_X1 U6905 ( .C1(n7486), .C2(n7430), .A(n7064), .B(n7063), .ZN(n7065)
         );
  OAI211_X1 U6906 ( .C1(alu_a_q[1]), .C2(alu_b_q[0]), .A(n7068), .B(alu_b_q[1]), .ZN(n7069) );
  OAI211_X1 U6907 ( .C1(n7774), .C2(n3804), .A(n7070), .B(n7069), .ZN(n7498)
         );
  INV_X1 U6908 ( .A(n7498), .ZN(n7380) );
  OAI222_X1 U6909 ( .A1(n3763), .A2(alu_a_q[2]), .B1(n3763), .B2(n7072), .C1(
        alu_a_q[2]), .C2(n7072), .ZN(n7096) );
  AOI22_X1 U6910 ( .A1(n3352), .A2(n7096), .B1(n3353), .B2(n7094), .ZN(n7075)
         );
  NAND2_X1 U6911 ( .A1(n3772), .A2(n3804), .ZN(n7095) );
  OAI22_X1 U6912 ( .A1(n7380), .A2(n7707), .B1(n7075), .B2(n7095), .ZN(n7092)
         );
  AOI22_X1 U6913 ( .A1(n3804), .A2(n7734), .B1(n7075), .B2(n7735), .ZN(n7076)
         );
  INV_X1 U6914 ( .A(n7076), .ZN(n7090) );
  NOR2_X1 U6915 ( .A1(n3794), .A2(n7883), .ZN(n7503) );
  NOR2_X1 U6916 ( .A1(n3785), .A2(n7774), .ZN(n7373) );
  NOR2_X1 U6917 ( .A1(n3786), .A2(n7122), .ZN(n7551) );
  NOR2_X1 U6918 ( .A1(n3793), .A2(n7082), .ZN(n7450) );
  NOR4_X1 U6919 ( .A1(n7503), .A2(n7373), .A3(n7551), .A4(n7450), .ZN(n7390)
         );
  INV_X1 U6920 ( .A(n7077), .ZN(n7877) );
  NAND2_X1 U6921 ( .A1(alu_a_q[13]), .A2(n7125), .ZN(n7375) );
  NAND2_X1 U6922 ( .A1(alu_a_q[11]), .A2(n7743), .ZN(n7264) );
  NAND2_X1 U6923 ( .A1(alu_a_q[14]), .A2(n7146), .ZN(n7447) );
  NAND2_X1 U6924 ( .A1(alu_a_q[12]), .A2(n7101), .ZN(n7309) );
  NAND4_X1 U6925 ( .A1(n7375), .A2(n7264), .A3(n7447), .A4(n7309), .ZN(n7263)
         );
  NAND2_X1 U6926 ( .A1(alu_a_q[9]), .A2(n7125), .ZN(n7267) );
  NAND2_X1 U6927 ( .A1(alu_a_q[7]), .A2(n7743), .ZN(n7171) );
  NAND2_X1 U6928 ( .A1(alu_a_q[8]), .A2(n7101), .ZN(n7214) );
  NAND2_X1 U6929 ( .A1(alu_a_q[10]), .A2(n7146), .ZN(n7308) );
  NAND4_X1 U6930 ( .A1(n7267), .A2(n7171), .A3(n7214), .A4(n7308), .ZN(n7168)
         );
  AOI22_X1 U6931 ( .A1(n7749), .A2(n7263), .B1(n7740), .B2(n7168), .ZN(n7080)
         );
  NOR2_X1 U6932 ( .A1(n3780), .A2(n7082), .ZN(n7124) );
  NAND2_X1 U6933 ( .A1(alu_a_q[5]), .A2(n7125), .ZN(n7169) );
  NAND2_X1 U6934 ( .A1(alu_a_q[6]), .A2(n7146), .ZN(n7217) );
  OAI211_X1 U6935 ( .C1(n7774), .C2(n3804), .A(n7169), .B(n7217), .ZN(n7078)
         );
  OAI21_X1 U6936 ( .B1(n7124), .B2(n7078), .A(n7748), .ZN(n7079) );
  OAI211_X1 U6937 ( .C1(n7390), .C2(n7877), .A(n7080), .B(n7079), .ZN(n7085)
         );
  NOR2_X1 U6938 ( .A1(n3766), .A2(n7883), .ZN(n7598) );
  NOR2_X1 U6939 ( .A1(n3787), .A2(n7774), .ZN(n7504) );
  NOR2_X1 U6940 ( .A1(n3795), .A2(n7122), .ZN(n7651) );
  NOR2_X1 U6941 ( .A1(n3791), .A2(n7082), .ZN(n7549) );
  NOR4_X1 U6942 ( .A1(n7598), .A2(n7504), .A3(n7651), .A4(n7549), .ZN(n7384)
         );
  NOR2_X1 U6943 ( .A1(n3831), .A2(n7774), .ZN(n7839) );
  OR2_X1 U6944 ( .A1(n7857), .A2(n7839), .ZN(n7387) );
  NOR2_X1 U6945 ( .A1(n3784), .A2(n7774), .ZN(n7705) );
  NOR2_X1 U6946 ( .A1(n3797), .A2(n7883), .ZN(n7837) );
  NOR2_X1 U6947 ( .A1(n3790), .A2(n7082), .ZN(n7776) );
  NOR2_X1 U6948 ( .A1(n3833), .A2(n7122), .ZN(n7081) );
  NOR4_X1 U6949 ( .A1(n7705), .A2(n7837), .A3(n7776), .A4(n7081), .ZN(n7382)
         );
  NOR2_X1 U6950 ( .A1(n3792), .A2(n7774), .ZN(n7597) );
  NOR2_X1 U6951 ( .A1(n3829), .A2(n7883), .ZN(n7706) );
  NOR2_X1 U6952 ( .A1(n3789), .A2(n7082), .ZN(n7650) );
  NOR2_X1 U6953 ( .A1(n3832), .A2(n7122), .ZN(n7775) );
  NOR4_X1 U6954 ( .A1(n7597), .A2(n7706), .A3(n7650), .A4(n7775), .ZN(n7392)
         );
  OAI22_X1 U6955 ( .A1(n7382), .A2(n7313), .B1(n7392), .B2(n7282), .ZN(n7083)
         );
  AOI21_X1 U6956 ( .B1(n7418), .B2(n7387), .A(n7083), .ZN(n7084) );
  OAI21_X1 U6957 ( .B1(n7384), .B2(n7427), .A(n7084), .ZN(n7511) );
  OAI221_X1 U6958 ( .B1(n7085), .B2(alu_b_q[4]), .C1(n7085), .C2(n7511), .A(
        n7887), .ZN(n7089) );
  OAI22_X1 U6959 ( .A1(n3764), .A2(n7096), .B1(n3842), .B2(n7094), .ZN(n7087)
         );
  NAND2_X1 U6960 ( .A1(alu_b_q[3]), .A2(alu_a_q[3]), .ZN(n7086) );
  OAI211_X1 U6961 ( .C1(n7835), .C2(n7087), .A(n7095), .B(n7086), .ZN(n7088)
         );
  OAI211_X1 U6962 ( .C1(n3772), .C2(n7090), .A(n7089), .B(n7088), .ZN(n7091)
         );
  NOR2_X1 U6963 ( .A1(alu_b_q[4]), .A2(alu_a_q[4]), .ZN(n7117) );
  OAI222_X1 U6964 ( .A1(n3804), .A2(n7096), .B1(n3804), .B2(alu_b_q[3]), .C1(
        n7096), .C2(alu_b_q[3]), .ZN(n7106) );
  OAI22_X1 U6965 ( .A1(n7116), .A2(n3842), .B1(n3764), .B2(n7106), .ZN(n7114)
         );
  NAND2_X1 U6966 ( .A1(alu_a_q[21]), .A2(n7101), .ZN(n7570) );
  NAND2_X1 U6967 ( .A1(alu_a_q[23]), .A2(n7146), .ZN(n7674) );
  NAND2_X1 U6968 ( .A1(alu_a_q[20]), .A2(n7743), .ZN(n7524) );
  NAND2_X1 U6969 ( .A1(alu_a_q[22]), .A2(n7125), .ZN(n7617) );
  NAND4_X1 U6970 ( .A1(n7570), .A2(n7674), .A3(n7524), .A4(n7617), .ZN(n7410)
         );
  NOR2_X1 U6971 ( .A1(n7429), .A2(n7379), .ZN(n7142) );
  NAND2_X1 U6972 ( .A1(alu_a_q[27]), .A2(n7146), .ZN(n7805) );
  NAND2_X1 U6973 ( .A1(alu_a_q[25]), .A2(n7101), .ZN(n7675) );
  NAND2_X1 U6974 ( .A1(alu_a_q[24]), .A2(n7743), .ZN(n7618) );
  NAND2_X1 U6975 ( .A1(alu_a_q[26]), .A2(n7125), .ZN(n7747) );
  NAND4_X1 U6976 ( .A1(n7805), .A2(n7675), .A3(n7618), .A4(n7747), .ZN(n7412)
         );
  INV_X1 U6977 ( .A(n7412), .ZN(n7284) );
  AOI22_X1 U6978 ( .A1(alu_a_q[30]), .A2(n7125), .B1(alu_a_q[31]), .B2(n7146), 
        .ZN(n7097) );
  NAND2_X1 U6979 ( .A1(alu_a_q[29]), .A2(n7101), .ZN(n7804) );
  OAI211_X1 U6980 ( .C1(n7774), .C2(n3790), .A(n7097), .B(n7804), .ZN(n7411)
         );
  INV_X1 U6981 ( .A(n7411), .ZN(n7197) );
  OAI22_X1 U6982 ( .A1(n7284), .A2(n7282), .B1(n7197), .B2(n7313), .ZN(n7098)
         );
  AOI211_X1 U6983 ( .C1(n7414), .C2(n7410), .A(n7142), .B(n7098), .ZN(n7529)
         );
  NOR2_X1 U6984 ( .A1(n3808), .A2(n7774), .ZN(n7428) );
  AOI22_X1 U6985 ( .A1(alu_a_q[3]), .A2(n7101), .B1(alu_a_q[1]), .B2(n7146), 
        .ZN(n7099) );
  NAND2_X1 U6986 ( .A1(alu_a_q[4]), .A2(n7743), .ZN(n7100) );
  OAI211_X1 U6987 ( .C1(n7883), .C2(n3803), .A(n7099), .B(n7100), .ZN(n7419)
         );
  AOI22_X1 U6988 ( .A1(alu_b_q[2]), .A2(n7428), .B1(n7419), .B2(n3763), .ZN(
        n7280) );
  NOR2_X1 U6989 ( .A1(alu_b_q[3]), .A2(n7280), .ZN(n7544) );
  NAND2_X1 U6990 ( .A1(alu_a_q[9]), .A2(n7101), .ZN(n7230) );
  NAND2_X1 U6991 ( .A1(alu_a_q[11]), .A2(n7146), .ZN(n7348) );
  NAND2_X1 U6992 ( .A1(alu_a_q[10]), .A2(n7125), .ZN(n7279) );
  NAND2_X1 U6993 ( .A1(alu_a_q[8]), .A2(n7743), .ZN(n7192) );
  AND4_X1 U6994 ( .A1(n7230), .A2(n7348), .A3(n7279), .A4(n7192), .ZN(n7880)
         );
  OAI22_X1 U6995 ( .A1(n7880), .A2(n7385), .B1(n3780), .B2(n7867), .ZN(n7104)
         );
  NAND2_X1 U6996 ( .A1(alu_a_q[15]), .A2(n7146), .ZN(n7476) );
  NAND2_X1 U6997 ( .A1(alu_a_q[13]), .A2(n7101), .ZN(n7347) );
  NAND2_X1 U6998 ( .A1(alu_a_q[12]), .A2(n7743), .ZN(n7278) );
  NAND2_X1 U6999 ( .A1(alu_a_q[14]), .A2(n7125), .ZN(n7422) );
  AND4_X1 U7000 ( .A1(n7476), .A2(n7347), .A3(n7278), .A4(n7422), .ZN(n7878)
         );
  INV_X1 U7001 ( .A(n7356), .ZN(n7391) );
  NAND2_X1 U7002 ( .A1(alu_a_q[5]), .A2(n7101), .ZN(n7149) );
  NAND2_X1 U7003 ( .A1(alu_a_q[7]), .A2(n7146), .ZN(n7231) );
  NAND2_X1 U7004 ( .A1(alu_a_q[6]), .A2(n7125), .ZN(n7191) );
  NAND4_X1 U7005 ( .A1(n7149), .A2(n7231), .A3(n7100), .A4(n7191), .ZN(n7873)
         );
  NAND2_X1 U7006 ( .A1(alu_a_q[19]), .A2(n7146), .ZN(n7571) );
  NAND2_X1 U7007 ( .A1(alu_a_q[17]), .A2(n7101), .ZN(n7477) );
  NAND2_X1 U7008 ( .A1(alu_a_q[16]), .A2(n7743), .ZN(n7423) );
  NAND2_X1 U7009 ( .A1(alu_a_q[18]), .A2(n7125), .ZN(n7525) );
  NAND4_X1 U7010 ( .A1(n7571), .A2(n7477), .A3(n7423), .A4(n7525), .ZN(n7413)
         );
  AOI22_X1 U7011 ( .A1(n7885), .A2(n7873), .B1(n7354), .B2(n7413), .ZN(n7102)
         );
  OAI21_X1 U7012 ( .B1(n7878), .B2(n7391), .A(n7102), .ZN(n7103) );
  AOI211_X1 U7013 ( .C1(n7425), .C2(n7544), .A(n7104), .B(n7103), .ZN(n7105)
         );
  OAI21_X1 U7014 ( .B1(n7529), .B2(n7430), .A(n7105), .ZN(n7113) );
  OAI21_X1 U7015 ( .B1(n7119), .B2(n3764), .A(n7865), .ZN(n7107) );
  AOI21_X1 U7016 ( .B1(n3353), .B2(n7116), .A(n7107), .ZN(n7111) );
  OR3_X1 U7017 ( .A1(n3780), .A2(n7114), .A3(n7342), .ZN(n7108) );
  NAND2_X1 U7018 ( .A1(n7108), .A2(alu_b_q[4]), .ZN(n7110) );
  NOR2_X1 U7019 ( .A1(alu_a_q[4]), .A2(n7872), .ZN(n7109) );
  NAND2_X1 U7020 ( .A1(alu_a_q[4]), .A2(n3809), .ZN(n7118) );
  AOI222_X1 U7021 ( .A1(n7111), .A2(n7110), .B1(n7111), .B2(n7109), .C1(n7110), 
        .C2(n7118), .ZN(n7112) );
  AOI21_X1 U7022 ( .B1(n3352), .B2(n7138), .A(n7835), .ZN(n7120) );
  OAI21_X1 U7023 ( .B1(n3842), .B2(n7140), .A(n7120), .ZN(n7136) );
  NAND2_X1 U7024 ( .A1(alu_b_q[5]), .A2(n3781), .ZN(n7139) );
  OAI21_X1 U7025 ( .B1(alu_b_q[5]), .B2(n3781), .A(n7139), .ZN(n7135) );
  INV_X1 U7026 ( .A(n7788), .ZN(n7871) );
  INV_X1 U7027 ( .A(n7138), .ZN(n7121) );
  AOI222_X1 U7028 ( .A1(n7140), .A2(n3353), .B1(alu_b_q[5]), .B2(n7871), .C1(
        n3352), .C2(n7121), .ZN(n7133) );
  OAI22_X1 U7029 ( .A1(n3781), .A2(n7774), .B1(n3803), .B2(n7122), .ZN(n7123)
         );
  AOI211_X1 U7030 ( .C1(n7125), .C2(alu_a_q[3]), .A(n7124), .B(n7123), .ZN(
        n7314) );
  INV_X1 U7031 ( .A(n7314), .ZN(n7452) );
  AOI22_X1 U7032 ( .A1(n7414), .A2(n7452), .B1(n7424), .B2(n7446), .ZN(n7547)
         );
  OAI22_X1 U7033 ( .A1(n7547), .A2(n7399), .B1(n7306), .B2(n7383), .ZN(n7131)
         );
  OAI22_X1 U7034 ( .A1(n7322), .A2(n7282), .B1(n7307), .B2(n7427), .ZN(n7126)
         );
  AOI211_X1 U7035 ( .C1(n7417), .C2(n7316), .A(n7142), .B(n7126), .ZN(n7554)
         );
  AOI22_X1 U7036 ( .A1(alu_b_q[5]), .A2(n7872), .B1(n7885), .B2(n7127), .ZN(
        n7129) );
  AOI22_X1 U7037 ( .A1(alu_a_q[5]), .A2(n7802), .B1(n7356), .B2(n7319), .ZN(
        n7128) );
  OAI211_X1 U7038 ( .C1(n7554), .C2(n7430), .A(n7129), .B(n7128), .ZN(n7130)
         );
  AOI211_X1 U7039 ( .C1(n7874), .C2(n7220), .A(n7131), .B(n7130), .ZN(n7132)
         );
  OAI21_X1 U7040 ( .B1(n7133), .B2(n7135), .A(n7132), .ZN(n7134) );
  NOR2_X1 U7041 ( .A1(alu_b_q[6]), .A2(n3773), .ZN(n7160) );
  OAI22_X1 U7042 ( .A1(n7162), .A2(n3764), .B1(n3842), .B2(n7164), .ZN(n7159)
         );
  AOI22_X1 U7043 ( .A1(n3352), .A2(n7162), .B1(n3353), .B2(n7164), .ZN(n7157)
         );
  NAND2_X1 U7044 ( .A1(n3773), .A2(n3810), .ZN(n7165) );
  INV_X1 U7045 ( .A(n7430), .ZN(n7947) );
  AOI22_X1 U7046 ( .A1(n7414), .A2(n7355), .B1(n7417), .B2(n7341), .ZN(n7144)
         );
  INV_X1 U7047 ( .A(n7142), .ZN(n7143) );
  OAI211_X1 U7048 ( .C1(n7352), .C2(n7282), .A(n7144), .B(n7143), .ZN(n7588)
         );
  AOI22_X1 U7049 ( .A1(n7874), .A2(n7234), .B1(n7356), .B2(n7358), .ZN(n7145)
         );
  OAI21_X1 U7050 ( .B1(n3773), .B2(n7867), .A(n7145), .ZN(n7153) );
  NAND2_X1 U7051 ( .A1(alu_a_q[3]), .A2(n7146), .ZN(n7882) );
  NAND4_X1 U7052 ( .A1(n7149), .A2(n7882), .A3(n7148), .A4(n7147), .ZN(n7479)
         );
  AOI22_X1 U7053 ( .A1(n7414), .A2(n7479), .B1(n7424), .B2(n7478), .ZN(n7573)
         );
  AOI22_X1 U7054 ( .A1(n7885), .A2(n7150), .B1(n7354), .B2(n7357), .ZN(n7151)
         );
  OAI21_X1 U7055 ( .B1(n7573), .B2(n7399), .A(n7151), .ZN(n7152) );
  AOI211_X1 U7056 ( .C1(n7947), .C2(n7588), .A(n7153), .B(n7152), .ZN(n7156)
         );
  NOR2_X1 U7057 ( .A1(alu_a_q[6]), .A2(n3810), .ZN(n7163) );
  AOI211_X1 U7058 ( .C1(n7735), .C2(n7157), .A(n3810), .B(n3773), .ZN(n7154)
         );
  AOI221_X1 U7059 ( .B1(n7624), .B2(n7163), .C1(n7159), .C2(n7163), .A(n7154), 
        .ZN(n7155) );
  OAI211_X1 U7060 ( .C1(n7157), .C2(n7165), .A(n7156), .B(n7155), .ZN(n7158)
         );
  AOI22_X1 U7061 ( .A1(n4847), .A2(n4828), .B1(n3876), .B2(n4846), .ZN(n2618)
         );
  AOI22_X1 U7062 ( .A1(n4849), .A2(n4828), .B1(n4396), .B2(n4848), .ZN(n2617)
         );
  AOI22_X1 U7063 ( .A1(n4851), .A2(n4828), .B1(n4184), .B2(n4850), .ZN(n2616)
         );
  AOI22_X1 U7064 ( .A1(n4853), .A2(n4828), .B1(n4185), .B2(n4852), .ZN(n2615)
         );
  AOI22_X1 U7065 ( .A1(n4855), .A2(n4828), .B1(n4397), .B2(n4854), .ZN(n2614)
         );
  AOI22_X1 U7066 ( .A1(n4857), .A2(n4828), .B1(n3877), .B2(n4856), .ZN(n2613)
         );
  AOI22_X1 U7067 ( .A1(n4859), .A2(n4828), .B1(n3878), .B2(n4858), .ZN(n2612)
         );
  AOI22_X1 U7068 ( .A1(n4861), .A2(n4828), .B1(n4398), .B2(n4860), .ZN(n2611)
         );
  AOI22_X1 U7069 ( .A1(n4863), .A2(n4828), .B1(n3879), .B2(n4862), .ZN(n2610)
         );
  AOI22_X1 U7070 ( .A1(n4865), .A2(n4828), .B1(n4399), .B2(n4864), .ZN(n2609)
         );
  AOI22_X1 U7071 ( .A1(n4867), .A2(n4828), .B1(n4186), .B2(n4866), .ZN(n2608)
         );
  AOI22_X1 U7072 ( .A1(n4869), .A2(n4828), .B1(n4187), .B2(n4868), .ZN(n2607)
         );
  AOI22_X1 U7073 ( .A1(n4871), .A2(n4828), .B1(n4400), .B2(n4870), .ZN(n2606)
         );
  AOI22_X1 U7074 ( .A1(n4873), .A2(n4828), .B1(n3880), .B2(n4872), .ZN(n2605)
         );
  AOI22_X1 U7075 ( .A1(n4875), .A2(n4828), .B1(n3881), .B2(n4874), .ZN(n2604)
         );
  AOI22_X1 U7076 ( .A1(n4877), .A2(n4828), .B1(n4401), .B2(n4876), .ZN(n2603)
         );
  AOI22_X1 U7077 ( .A1(n4879), .A2(n4828), .B1(n3882), .B2(n4878), .ZN(n2602)
         );
  AOI22_X1 U7078 ( .A1(n4881), .A2(n4828), .B1(n4402), .B2(n4880), .ZN(n2601)
         );
  AOI22_X1 U7079 ( .A1(n4883), .A2(n4828), .B1(n4188), .B2(n4882), .ZN(n2600)
         );
  AOI22_X1 U7080 ( .A1(n4885), .A2(n4828), .B1(n4189), .B2(n4884), .ZN(n2599)
         );
  AOI22_X1 U7081 ( .A1(n4887), .A2(n4828), .B1(n4403), .B2(n4886), .ZN(n2598)
         );
  AOI22_X1 U7082 ( .A1(n4889), .A2(n7161), .B1(n3883), .B2(n4888), .ZN(n2597)
         );
  AOI22_X1 U7083 ( .A1(n4891), .A2(n7161), .B1(n3884), .B2(n4890), .ZN(n2596)
         );
  AOI22_X1 U7084 ( .A1(n4893), .A2(n7161), .B1(n4404), .B2(n4892), .ZN(n2595)
         );
  AOI22_X1 U7085 ( .A1(n7978), .A2(n7161), .B1(n3885), .B2(n4894), .ZN(n2594)
         );
  AOI22_X1 U7086 ( .A1(n7979), .A2(n7161), .B1(n4405), .B2(n4896), .ZN(n2593)
         );
  AOI22_X1 U7087 ( .A1(n7980), .A2(n7161), .B1(n4190), .B2(n4898), .ZN(n2592)
         );
  AOI22_X1 U7088 ( .A1(n7981), .A2(n4828), .B1(n4191), .B2(n4900), .ZN(n2591)
         );
  AOI22_X1 U7089 ( .A1(n7982), .A2(n4828), .B1(n4406), .B2(n4902), .ZN(n2590)
         );
  AOI22_X1 U7090 ( .A1(n7983), .A2(n4828), .B1(n3886), .B2(n4904), .ZN(n2589)
         );
  AOI22_X1 U7091 ( .A1(n7984), .A2(n4828), .B1(n3887), .B2(n4906), .ZN(n2588)
         );
  AOI22_X1 U7092 ( .A1(n7985), .A2(n4828), .B1(n4407), .B2(n4908), .ZN(n2587)
         );
  AOI22_X1 U7093 ( .A1(n3352), .A2(n7185), .B1(n3353), .B2(n7187), .ZN(n7166)
         );
  NOR2_X1 U7094 ( .A1(alu_a_q[7]), .A2(alu_b_q[7]), .ZN(n7188) );
  AOI21_X1 U7095 ( .B1(n7166), .B2(n7865), .A(n7188), .ZN(n7183) );
  NAND2_X1 U7096 ( .A1(alu_a_q[7]), .A2(alu_b_q[7]), .ZN(n7186) );
  NOR2_X1 U7097 ( .A1(n3772), .A2(n7429), .ZN(n7261) );
  OAI22_X1 U7098 ( .A1(n7382), .A2(n7282), .B1(n7392), .B2(n7427), .ZN(n7167)
         );
  AOI211_X1 U7099 ( .C1(n7839), .C2(n7417), .A(n7261), .B(n7167), .ZN(n7606)
         );
  NOR2_X1 U7100 ( .A1(n7380), .A2(n7282), .ZN(n7604) );
  AOI22_X1 U7101 ( .A1(n7425), .A2(n7604), .B1(n7885), .B2(n7168), .ZN(n7177)
         );
  OAI22_X1 U7102 ( .A1(n7384), .A2(n7383), .B1(n7390), .B2(n7391), .ZN(n7175)
         );
  NAND4_X1 U7103 ( .A1(n7172), .A2(n7171), .A3(n7170), .A4(n7169), .ZN(n7596)
         );
  INV_X1 U7104 ( .A(n7596), .ZN(n7500) );
  AOI22_X1 U7105 ( .A1(alu_b_q[7]), .A2(n7872), .B1(n7874), .B2(n7263), .ZN(
        n7173) );
  OAI21_X1 U7106 ( .B1(n7500), .B2(n7707), .A(n7173), .ZN(n7174) );
  AOI211_X1 U7107 ( .C1(alu_a_q[7]), .C2(n7802), .A(n7175), .B(n7174), .ZN(
        n7176) );
  OAI211_X1 U7108 ( .C1(n7606), .C2(n7430), .A(n7177), .B(n7176), .ZN(n7182)
         );
  OAI22_X1 U7109 ( .A1(n3764), .A2(n7185), .B1(n3842), .B2(n7187), .ZN(n7179)
         );
  INV_X1 U7110 ( .A(n7186), .ZN(n7178) );
  OAI222_X1 U7111 ( .A1(n7179), .A2(n7178), .B1(n7179), .B2(n7871), .C1(n7178), 
        .C2(n7188), .ZN(n7180) );
  INV_X1 U7112 ( .A(n7180), .ZN(n7181) );
  AOI22_X1 U7113 ( .A1(n4847), .A2(n4829), .B1(n3888), .B2(n4846), .ZN(n2586)
         );
  AOI22_X1 U7114 ( .A1(n4849), .A2(n4829), .B1(n4408), .B2(n4848), .ZN(n2585)
         );
  AOI22_X1 U7115 ( .A1(n4851), .A2(n4829), .B1(n4192), .B2(n4850), .ZN(n2584)
         );
  AOI22_X1 U7116 ( .A1(n4853), .A2(n4829), .B1(n4193), .B2(n4852), .ZN(n2583)
         );
  AOI22_X1 U7117 ( .A1(n4855), .A2(n4829), .B1(n4409), .B2(n4854), .ZN(n2582)
         );
  AOI22_X1 U7118 ( .A1(n4857), .A2(n4829), .B1(n3889), .B2(n4856), .ZN(n2581)
         );
  AOI22_X1 U7119 ( .A1(n4859), .A2(n4829), .B1(n3890), .B2(n4858), .ZN(n2580)
         );
  AOI22_X1 U7120 ( .A1(n4861), .A2(n4829), .B1(n4410), .B2(n4860), .ZN(n2579)
         );
  AOI22_X1 U7121 ( .A1(n4863), .A2(n4829), .B1(n3891), .B2(n4862), .ZN(n2578)
         );
  AOI22_X1 U7122 ( .A1(n4865), .A2(n4829), .B1(n4411), .B2(n4864), .ZN(n2577)
         );
  AOI22_X1 U7123 ( .A1(n4867), .A2(n4829), .B1(n4194), .B2(n4866), .ZN(n2576)
         );
  AOI22_X1 U7124 ( .A1(n4869), .A2(n4829), .B1(n4195), .B2(n4868), .ZN(n2575)
         );
  AOI22_X1 U7125 ( .A1(n4871), .A2(n4829), .B1(n4412), .B2(n4870), .ZN(n2574)
         );
  AOI22_X1 U7126 ( .A1(n4873), .A2(n4829), .B1(n3892), .B2(n4872), .ZN(n2573)
         );
  AOI22_X1 U7127 ( .A1(n4875), .A2(n4829), .B1(n3893), .B2(n4874), .ZN(n2572)
         );
  AOI22_X1 U7128 ( .A1(n4877), .A2(n4829), .B1(n4413), .B2(n4876), .ZN(n2571)
         );
  AOI22_X1 U7129 ( .A1(n7970), .A2(n4829), .B1(n3894), .B2(n4878), .ZN(n2570)
         );
  AOI22_X1 U7130 ( .A1(n7971), .A2(n4829), .B1(n4414), .B2(n4880), .ZN(n2569)
         );
  AOI22_X1 U7131 ( .A1(n7972), .A2(n4829), .B1(n4196), .B2(n4882), .ZN(n2568)
         );
  AOI22_X1 U7132 ( .A1(n7973), .A2(n4829), .B1(n4197), .B2(n4884), .ZN(n2567)
         );
  AOI22_X1 U7133 ( .A1(n7974), .A2(n4829), .B1(n4415), .B2(n4886), .ZN(n2566)
         );
  AOI22_X1 U7134 ( .A1(n7975), .A2(n7184), .B1(n3895), .B2(n4888), .ZN(n2565)
         );
  AOI22_X1 U7135 ( .A1(n7976), .A2(n7184), .B1(n3896), .B2(n4890), .ZN(n2564)
         );
  AOI22_X1 U7136 ( .A1(n7977), .A2(n7184), .B1(n4416), .B2(n4892), .ZN(n2563)
         );
  AOI22_X1 U7137 ( .A1(n7978), .A2(n7184), .B1(n3897), .B2(n4894), .ZN(n2562)
         );
  AOI22_X1 U7138 ( .A1(n7979), .A2(n7184), .B1(n4417), .B2(n4896), .ZN(n2561)
         );
  AOI22_X1 U7139 ( .A1(n7980), .A2(n7184), .B1(n4198), .B2(n4898), .ZN(n2560)
         );
  AOI22_X1 U7140 ( .A1(n7981), .A2(n4829), .B1(n4199), .B2(n4900), .ZN(n2559)
         );
  AOI22_X1 U7141 ( .A1(n7982), .A2(n4829), .B1(n4418), .B2(n4902), .ZN(n2558)
         );
  AOI22_X1 U7142 ( .A1(n7983), .A2(n4829), .B1(n3898), .B2(n4904), .ZN(n2557)
         );
  AOI22_X1 U7143 ( .A1(n7984), .A2(n4829), .B1(n3899), .B2(n4906), .ZN(n2556)
         );
  AOI22_X1 U7144 ( .A1(n7985), .A2(n4829), .B1(n4419), .B2(n4908), .ZN(n2555)
         );
  AOI222_X1 U7145 ( .A1(alu_a_q[7]), .A2(n3814), .B1(alu_a_q[7]), .B2(n7185), 
        .C1(n3814), .C2(n7185), .ZN(n7210) );
  AOI22_X1 U7146 ( .A1(n3352), .A2(n7210), .B1(n3353), .B2(n7208), .ZN(n7199)
         );
  AOI211_X1 U7147 ( .C1(n7735), .C2(n7199), .A(n3805), .B(n3778), .ZN(n7206)
         );
  NAND4_X1 U7148 ( .A1(n7192), .A2(n7191), .A3(n7190), .A4(n7189), .ZN(n7521)
         );
  AOI222_X1 U7149 ( .A1(n7521), .A2(n7414), .B1(n7417), .B2(n7428), .C1(n7419), 
        .C2(n7424), .ZN(n7633) );
  INV_X1 U7150 ( .A(n7413), .ZN(n7193) );
  OAI22_X1 U7151 ( .A1(n7193), .A2(n7391), .B1(n7880), .B2(n7389), .ZN(n7195)
         );
  OAI22_X1 U7152 ( .A1(n7878), .A2(n7385), .B1(n3778), .B2(n7867), .ZN(n7194)
         );
  AOI211_X1 U7153 ( .C1(n7354), .C2(n7410), .A(n7195), .B(n7194), .ZN(n7196)
         );
  OAI21_X1 U7154 ( .B1(n7633), .B2(n7399), .A(n7196), .ZN(n7205) );
  INV_X1 U7155 ( .A(n7261), .ZN(n7232) );
  OAI21_X1 U7156 ( .B1(n7197), .B2(n7282), .A(n7232), .ZN(n7198) );
  AOI21_X1 U7157 ( .B1(n7414), .B2(n7412), .A(n7198), .ZN(n7632) );
  NAND2_X1 U7158 ( .A1(n3778), .A2(n3805), .ZN(n7209) );
  OAI22_X1 U7159 ( .A1(n7632), .A2(n7430), .B1(n7199), .B2(n7209), .ZN(n7204)
         );
  OAI22_X1 U7160 ( .A1(n7210), .A2(n3764), .B1(n3842), .B2(n7208), .ZN(n7200)
         );
  NOR2_X1 U7161 ( .A1(alu_a_q[8]), .A2(n3805), .ZN(n7211) );
  OAI21_X1 U7162 ( .B1(n7200), .B2(n7624), .A(n7211), .ZN(n7202) );
  OAI211_X1 U7163 ( .C1(n7835), .C2(n7200), .A(alu_a_q[8]), .B(n3805), .ZN(
        n7201) );
  NAND2_X1 U7164 ( .A1(n7202), .A2(n7201), .ZN(n7203) );
  NOR4_X1 U7165 ( .A1(n7206), .A2(n7205), .A3(n7204), .A4(n7203), .ZN(n7207)
         );
  AOI22_X1 U7166 ( .A1(n7954), .A2(n3370), .B1(n3900), .B2(n4846), .ZN(n2554)
         );
  AOI22_X1 U7167 ( .A1(n7955), .A2(n3370), .B1(n4420), .B2(n4848), .ZN(n2553)
         );
  AOI22_X1 U7168 ( .A1(n7956), .A2(n3370), .B1(n4200), .B2(n4850), .ZN(n2552)
         );
  AOI22_X1 U7169 ( .A1(n7957), .A2(n3370), .B1(n4201), .B2(n4852), .ZN(n2551)
         );
  AOI22_X1 U7170 ( .A1(n7958), .A2(n3370), .B1(n4421), .B2(n4854), .ZN(n2550)
         );
  AOI22_X1 U7171 ( .A1(n7959), .A2(n3370), .B1(n3901), .B2(n4856), .ZN(n2549)
         );
  AOI22_X1 U7172 ( .A1(n7960), .A2(n3370), .B1(n3902), .B2(n4858), .ZN(n2548)
         );
  AOI22_X1 U7173 ( .A1(n7961), .A2(n3370), .B1(n4422), .B2(n4860), .ZN(n2547)
         );
  AOI22_X1 U7174 ( .A1(n7962), .A2(n3370), .B1(n3903), .B2(n4862), .ZN(n2546)
         );
  AOI22_X1 U7175 ( .A1(n7963), .A2(n3370), .B1(n4423), .B2(n4864), .ZN(n2545)
         );
  AOI22_X1 U7176 ( .A1(n7964), .A2(n3370), .B1(n4202), .B2(n4866), .ZN(n2544)
         );
  AOI22_X1 U7177 ( .A1(n7965), .A2(n3370), .B1(n4203), .B2(n4868), .ZN(n2543)
         );
  AOI22_X1 U7178 ( .A1(n7966), .A2(n7207), .B1(n4424), .B2(n4870), .ZN(n2542)
         );
  AOI22_X1 U7179 ( .A1(n7967), .A2(n3370), .B1(n3904), .B2(n4872), .ZN(n2541)
         );
  AOI22_X1 U7180 ( .A1(n7968), .A2(n3370), .B1(n3905), .B2(n4874), .ZN(n2540)
         );
  AOI22_X1 U7181 ( .A1(n7969), .A2(n3370), .B1(n4425), .B2(n4876), .ZN(n2539)
         );
  AOI22_X1 U7182 ( .A1(n7970), .A2(n3370), .B1(n3906), .B2(n4878), .ZN(n2538)
         );
  AOI22_X1 U7183 ( .A1(n7971), .A2(n3370), .B1(n4426), .B2(n4880), .ZN(n2537)
         );
  AOI22_X1 U7184 ( .A1(n7972), .A2(n3370), .B1(n4204), .B2(n4882), .ZN(n2536)
         );
  AOI22_X1 U7185 ( .A1(n7973), .A2(n3370), .B1(n4205), .B2(n4884), .ZN(n2535)
         );
  AOI22_X1 U7186 ( .A1(n7974), .A2(n3370), .B1(n4427), .B2(n4886), .ZN(n2534)
         );
  AOI22_X1 U7187 ( .A1(n7975), .A2(n3370), .B1(n3907), .B2(n4888), .ZN(n2533)
         );
  AOI22_X1 U7188 ( .A1(n7976), .A2(n3370), .B1(n3908), .B2(n4890), .ZN(n2532)
         );
  AOI22_X1 U7189 ( .A1(n7977), .A2(n3370), .B1(n4428), .B2(n4892), .ZN(n2531)
         );
  AOI22_X1 U7190 ( .A1(n7978), .A2(n3370), .B1(n3909), .B2(n4894), .ZN(n2530)
         );
  AOI22_X1 U7191 ( .A1(n7979), .A2(n3370), .B1(n4429), .B2(n4896), .ZN(n2529)
         );
  AOI22_X1 U7192 ( .A1(n7980), .A2(n3370), .B1(n4206), .B2(n4898), .ZN(n2528)
         );
  AOI22_X1 U7193 ( .A1(n4901), .A2(n3370), .B1(n4207), .B2(n4900), .ZN(n2527)
         );
  AOI22_X1 U7194 ( .A1(n4903), .A2(n3370), .B1(n4430), .B2(n4902), .ZN(n2526)
         );
  AOI22_X1 U7195 ( .A1(n7983), .A2(n3370), .B1(n3910), .B2(n4904), .ZN(n2525)
         );
  AOI22_X1 U7196 ( .A1(n4907), .A2(n3370), .B1(n3911), .B2(n4906), .ZN(n2524)
         );
  AOI22_X1 U7197 ( .A1(n7985), .A2(n3370), .B1(n4431), .B2(n4908), .ZN(n2523)
         );
  NOR2_X1 U7198 ( .A1(alu_a_q[9]), .A2(alu_b_q[9]), .ZN(n7242) );
  OAI22_X1 U7199 ( .A1(alu_b_q[8]), .A2(n3778), .B1(n7211), .B2(n7210), .ZN(
        n7238) );
  OAI22_X1 U7200 ( .A1(n7241), .A2(n3842), .B1(n3764), .B2(n7238), .ZN(n7226)
         );
  AOI22_X1 U7201 ( .A1(n3352), .A2(n7238), .B1(n3353), .B2(n7241), .ZN(n7212)
         );
  NAND2_X1 U7202 ( .A1(n3782), .A2(alu_a_q[9]), .ZN(n7240) );
  AOI21_X1 U7203 ( .B1(n7212), .B2(n7865), .A(n7240), .ZN(n7225) );
  INV_X1 U7204 ( .A(n7624), .ZN(n7676) );
  AOI22_X1 U7205 ( .A1(alu_a_q[9]), .A2(n7802), .B1(n7874), .B2(n7319), .ZN(
        n7222) );
  OAI22_X1 U7206 ( .A1(n7306), .A2(n7391), .B1(n7307), .B2(n7383), .ZN(n7219)
         );
  OAI21_X1 U7207 ( .B1(n7322), .B2(n7427), .A(n7232), .ZN(n7213) );
  AOI21_X1 U7208 ( .B1(n7424), .B2(n7316), .A(n7213), .ZN(n7647) );
  NAND4_X1 U7209 ( .A1(n7217), .A2(n7216), .A3(n7215), .A4(n7214), .ZN(n7552)
         );
  AOI222_X1 U7210 ( .A1(n7552), .A2(n7414), .B1(n7446), .B2(n7417), .C1(n7452), 
        .C2(n7424), .ZN(n7646) );
  OAI22_X1 U7211 ( .A1(n7647), .A2(n7430), .B1(n7646), .B2(n7399), .ZN(n7218)
         );
  AOI211_X1 U7212 ( .C1(n7885), .C2(n7220), .A(n7219), .B(n7218), .ZN(n7221)
         );
  OAI211_X1 U7213 ( .C1(n3782), .C2(n7223), .A(n7222), .B(n7221), .ZN(n7224)
         );
  AOI22_X1 U7214 ( .A1(n7954), .A2(n4830), .B1(n3912), .B2(n4846), .ZN(n2522)
         );
  AOI22_X1 U7215 ( .A1(n7955), .A2(n4830), .B1(n4432), .B2(n4848), .ZN(n2521)
         );
  AOI22_X1 U7216 ( .A1(n7956), .A2(n4830), .B1(n4208), .B2(n4850), .ZN(n2520)
         );
  AOI22_X1 U7217 ( .A1(n7957), .A2(n4830), .B1(n4209), .B2(n4852), .ZN(n2519)
         );
  AOI22_X1 U7218 ( .A1(n7958), .A2(n4830), .B1(n4433), .B2(n4854), .ZN(n2518)
         );
  AOI22_X1 U7219 ( .A1(n7959), .A2(n4830), .B1(n3913), .B2(n4856), .ZN(n2517)
         );
  AOI22_X1 U7220 ( .A1(n7960), .A2(n4830), .B1(n3914), .B2(n4858), .ZN(n2516)
         );
  AOI22_X1 U7221 ( .A1(n7961), .A2(n4830), .B1(n4434), .B2(n4860), .ZN(n2515)
         );
  AOI22_X1 U7222 ( .A1(n7962), .A2(n4830), .B1(n3915), .B2(n4862), .ZN(n2514)
         );
  AOI22_X1 U7223 ( .A1(n7963), .A2(n4830), .B1(n4435), .B2(n4864), .ZN(n2513)
         );
  AOI22_X1 U7224 ( .A1(n7964), .A2(n4830), .B1(n4210), .B2(n4866), .ZN(n2512)
         );
  AOI22_X1 U7225 ( .A1(n7965), .A2(n4830), .B1(n4211), .B2(n4868), .ZN(n2511)
         );
  AOI22_X1 U7226 ( .A1(n7966), .A2(n4830), .B1(n4436), .B2(n4870), .ZN(n2510)
         );
  AOI22_X1 U7227 ( .A1(n7967), .A2(n4830), .B1(n3916), .B2(n4872), .ZN(n2509)
         );
  AOI22_X1 U7228 ( .A1(n7968), .A2(n4830), .B1(n3917), .B2(n4874), .ZN(n2508)
         );
  AOI22_X1 U7229 ( .A1(n7969), .A2(n4830), .B1(n4437), .B2(n4876), .ZN(n2507)
         );
  AOI22_X1 U7230 ( .A1(n7970), .A2(n4830), .B1(n3918), .B2(n4878), .ZN(n2506)
         );
  AOI22_X1 U7231 ( .A1(n7971), .A2(n4830), .B1(n4438), .B2(n4880), .ZN(n2505)
         );
  AOI22_X1 U7232 ( .A1(n7972), .A2(n4830), .B1(n4212), .B2(n4882), .ZN(n2504)
         );
  AOI22_X1 U7233 ( .A1(n7973), .A2(n4830), .B1(n4213), .B2(n4884), .ZN(n2503)
         );
  AOI22_X1 U7234 ( .A1(n7974), .A2(n4830), .B1(n4439), .B2(n4886), .ZN(n2502)
         );
  AOI22_X1 U7235 ( .A1(n7975), .A2(n7227), .B1(n3919), .B2(n4888), .ZN(n2501)
         );
  AOI22_X1 U7236 ( .A1(n7976), .A2(n7227), .B1(n3920), .B2(n4890), .ZN(n2500)
         );
  AOI22_X1 U7237 ( .A1(n7977), .A2(n7227), .B1(n4440), .B2(n4892), .ZN(n2499)
         );
  AOI22_X1 U7238 ( .A1(n7978), .A2(n7227), .B1(n3921), .B2(n4894), .ZN(n2498)
         );
  AOI22_X1 U7239 ( .A1(n7979), .A2(n7227), .B1(n4441), .B2(n4896), .ZN(n2497)
         );
  AOI22_X1 U7240 ( .A1(n7980), .A2(n7227), .B1(n4214), .B2(n4898), .ZN(n2496)
         );
  AOI22_X1 U7241 ( .A1(n4901), .A2(n4830), .B1(n4215), .B2(n4900), .ZN(n2495)
         );
  AOI22_X1 U7242 ( .A1(n4903), .A2(n4830), .B1(n4442), .B2(n4902), .ZN(n2494)
         );
  AOI22_X1 U7243 ( .A1(n4905), .A2(n4830), .B1(n3922), .B2(n4904), .ZN(n2493)
         );
  AOI22_X1 U7244 ( .A1(n4907), .A2(n4830), .B1(n3923), .B2(n4906), .ZN(n2492)
         );
  AOI22_X1 U7245 ( .A1(n4909), .A2(n4830), .B1(n4443), .B2(n4908), .ZN(n2491)
         );
  NAND4_X1 U7246 ( .A1(n7231), .A2(n7230), .A3(n7229), .A4(n7228), .ZN(n7581)
         );
  AOI222_X1 U7247 ( .A1(n7581), .A2(n7414), .B1(n7478), .B2(n7417), .C1(n7479), 
        .C2(n7424), .ZN(n7684) );
  OAI21_X1 U7248 ( .B1(n7352), .B2(n7427), .A(n7232), .ZN(n7233) );
  AOI21_X1 U7249 ( .B1(n7424), .B2(n7341), .A(n7233), .ZN(n7683) );
  OAI22_X1 U7250 ( .A1(n7684), .A2(n7399), .B1(n7683), .B2(n7430), .ZN(n7250)
         );
  AOI22_X1 U7251 ( .A1(alu_a_q[10]), .A2(n7802), .B1(alu_b_q[10]), .B2(n7872), 
        .ZN(n7237) );
  AOI22_X1 U7252 ( .A1(n7885), .A2(n7234), .B1(n7356), .B2(n7357), .ZN(n7236)
         );
  AOI22_X1 U7253 ( .A1(n7874), .A2(n7358), .B1(n7354), .B2(n7355), .ZN(n7235)
         );
  NAND3_X1 U7254 ( .A1(n7237), .A2(n7236), .A3(n7235), .ZN(n7249) );
  INV_X1 U7255 ( .A(n7238), .ZN(n7239) );
  INV_X1 U7256 ( .A(n7899), .ZN(n7243) );
  AOI222_X1 U7257 ( .A1(n7243), .A2(n3352), .B1(alu_a_q[10]), .B2(n7871), .C1(
        n7252), .C2(n3353), .ZN(n7247) );
  NAND2_X1 U7258 ( .A1(alu_a_q[10]), .A2(n3844), .ZN(n7290) );
  NOR2_X1 U7259 ( .A1(alu_a_q[10]), .A2(n3844), .ZN(n7893) );
  INV_X1 U7260 ( .A(n7893), .ZN(n7253) );
  NAND2_X1 U7261 ( .A1(n7290), .A2(n7253), .ZN(n7246) );
  OAI22_X1 U7262 ( .A1(n3764), .A2(n7243), .B1(n3842), .B2(n7252), .ZN(n7244)
         );
  OAI21_X1 U7263 ( .B1(n7244), .B2(n7835), .A(n7246), .ZN(n7245) );
  OAI21_X1 U7264 ( .B1(n7247), .B2(n7246), .A(n7245), .ZN(n7248) );
  AOI22_X1 U7265 ( .A1(n7954), .A2(n4831), .B1(n3924), .B2(n4846), .ZN(n2490)
         );
  AOI22_X1 U7266 ( .A1(n7955), .A2(n4831), .B1(n4444), .B2(n4848), .ZN(n2489)
         );
  AOI22_X1 U7267 ( .A1(n7956), .A2(n4831), .B1(n4216), .B2(n4850), .ZN(n2488)
         );
  AOI22_X1 U7268 ( .A1(n7957), .A2(n4831), .B1(n4217), .B2(n4852), .ZN(n2487)
         );
  AOI22_X1 U7269 ( .A1(n7958), .A2(n4831), .B1(n4445), .B2(n4854), .ZN(n2486)
         );
  AOI22_X1 U7270 ( .A1(n7959), .A2(n4831), .B1(n3925), .B2(n4856), .ZN(n2485)
         );
  AOI22_X1 U7271 ( .A1(n7960), .A2(n4831), .B1(n3926), .B2(n4858), .ZN(n2484)
         );
  AOI22_X1 U7272 ( .A1(n7961), .A2(n4831), .B1(n4446), .B2(n4860), .ZN(n2483)
         );
  AOI22_X1 U7273 ( .A1(n7962), .A2(n4831), .B1(n3927), .B2(n4862), .ZN(n2482)
         );
  AOI22_X1 U7274 ( .A1(n7963), .A2(n4831), .B1(n4447), .B2(n4864), .ZN(n2481)
         );
  AOI22_X1 U7275 ( .A1(n7964), .A2(n4831), .B1(n4218), .B2(n4866), .ZN(n2480)
         );
  AOI22_X1 U7276 ( .A1(n7965), .A2(n4831), .B1(n4219), .B2(n4868), .ZN(n2479)
         );
  AOI22_X1 U7277 ( .A1(n7966), .A2(n4831), .B1(n4448), .B2(n4870), .ZN(n2478)
         );
  AOI22_X1 U7278 ( .A1(n7967), .A2(n4831), .B1(n3928), .B2(n4872), .ZN(n2477)
         );
  AOI22_X1 U7279 ( .A1(n7968), .A2(n4831), .B1(n3929), .B2(n4874), .ZN(n2476)
         );
  AOI22_X1 U7280 ( .A1(n7969), .A2(n4831), .B1(n4449), .B2(n4876), .ZN(n2475)
         );
  AOI22_X1 U7281 ( .A1(n7970), .A2(n4831), .B1(n3930), .B2(n4878), .ZN(n2474)
         );
  AOI22_X1 U7282 ( .A1(n7971), .A2(n4831), .B1(n4450), .B2(n4880), .ZN(n2473)
         );
  AOI22_X1 U7283 ( .A1(n7972), .A2(n4831), .B1(n4220), .B2(n4882), .ZN(n2472)
         );
  AOI22_X1 U7284 ( .A1(n7973), .A2(n4831), .B1(n4221), .B2(n4884), .ZN(n2471)
         );
  AOI22_X1 U7285 ( .A1(n7974), .A2(n7251), .B1(n4451), .B2(n4886), .ZN(n2470)
         );
  AOI22_X1 U7286 ( .A1(n7975), .A2(n7251), .B1(n3931), .B2(n4888), .ZN(n2469)
         );
  AOI22_X1 U7287 ( .A1(n7976), .A2(n7251), .B1(n3932), .B2(n4890), .ZN(n2468)
         );
  AOI22_X1 U7288 ( .A1(n7977), .A2(n7251), .B1(n4452), .B2(n4892), .ZN(n2467)
         );
  AOI22_X1 U7289 ( .A1(n7978), .A2(n7251), .B1(n3933), .B2(n4894), .ZN(n2466)
         );
  AOI22_X1 U7290 ( .A1(n7979), .A2(n7251), .B1(n4453), .B2(n4896), .ZN(n2465)
         );
  AOI22_X1 U7291 ( .A1(n7980), .A2(n7251), .B1(n4222), .B2(n4898), .ZN(n2464)
         );
  AOI22_X1 U7292 ( .A1(n7981), .A2(n4831), .B1(n4223), .B2(n4900), .ZN(n2463)
         );
  AOI22_X1 U7293 ( .A1(n7982), .A2(n4831), .B1(n4454), .B2(n4902), .ZN(n2462)
         );
  AOI22_X1 U7294 ( .A1(n7983), .A2(n4831), .B1(n3934), .B2(n4904), .ZN(n2461)
         );
  AOI22_X1 U7295 ( .A1(n7984), .A2(n4831), .B1(n3935), .B2(n4906), .ZN(n2460)
         );
  AOI22_X1 U7296 ( .A1(n7985), .A2(n4831), .B1(n4455), .B2(n4908), .ZN(n2459)
         );
  NOR2_X1 U7297 ( .A1(alu_a_q[11]), .A2(alu_b_q[11]), .ZN(n7292) );
  NAND2_X1 U7298 ( .A1(n7290), .A2(n7289), .ZN(n7254) );
  OAI22_X1 U7299 ( .A1(n7293), .A2(n3842), .B1(n3764), .B2(n7254), .ZN(n7274)
         );
  AOI21_X1 U7300 ( .B1(n7254), .B2(n3352), .A(n7835), .ZN(n7255) );
  INV_X1 U7301 ( .A(n7255), .ZN(n7256) );
  AOI21_X1 U7302 ( .B1(n3353), .B2(n7293), .A(n7256), .ZN(n7260) );
  NAND2_X1 U7303 ( .A1(alu_a_q[11]), .A2(n7735), .ZN(n7257) );
  OAI21_X1 U7304 ( .B1(n7274), .B2(n7257), .A(alu_b_q[11]), .ZN(n7259) );
  NOR2_X1 U7305 ( .A1(alu_a_q[11]), .A2(n7872), .ZN(n7258) );
  NAND2_X1 U7306 ( .A1(alu_a_q[11]), .A2(n3775), .ZN(n7892) );
  AOI222_X1 U7307 ( .A1(n7260), .A2(n7259), .B1(n7260), .B2(n7258), .C1(n7259), 
        .C2(n7892), .ZN(n7273) );
  OAI21_X1 U7308 ( .B1(n7424), .B2(n7261), .A(n7387), .ZN(n7262) );
  OAI21_X1 U7309 ( .B1(n7382), .B2(n7427), .A(n7262), .ZN(n7698) );
  AOI22_X1 U7310 ( .A1(n7947), .A2(n7698), .B1(n7885), .B2(n7263), .ZN(n7271)
         );
  OAI22_X1 U7311 ( .A1(n7380), .A2(n7313), .B1(n7500), .B2(n7282), .ZN(n7697)
         );
  NAND4_X1 U7312 ( .A1(n7267), .A2(n7266), .A3(n7265), .A4(n7264), .ZN(n7700)
         );
  INV_X1 U7313 ( .A(n7700), .ZN(n7505) );
  OAI22_X1 U7314 ( .A1(n7505), .A2(n7707), .B1(n7392), .B2(n7383), .ZN(n7269)
         );
  OAI22_X1 U7315 ( .A1(n7390), .A2(n7385), .B1(n3813), .B2(n7867), .ZN(n7268)
         );
  AOI211_X1 U7316 ( .C1(n7425), .C2(n7697), .A(n7269), .B(n7268), .ZN(n7270)
         );
  OAI211_X1 U7317 ( .C1(n7384), .C2(n7391), .A(n7271), .B(n7270), .ZN(n7272)
         );
  AOI22_X1 U7318 ( .A1(n4847), .A2(n4832), .B1(n3936), .B2(n4846), .ZN(n2458)
         );
  AOI22_X1 U7319 ( .A1(n4849), .A2(n4832), .B1(n4456), .B2(n4848), .ZN(n2457)
         );
  AOI22_X1 U7320 ( .A1(n4851), .A2(n4832), .B1(n4224), .B2(n4850), .ZN(n2456)
         );
  AOI22_X1 U7321 ( .A1(n4853), .A2(n4832), .B1(n4225), .B2(n4852), .ZN(n2455)
         );
  AOI22_X1 U7322 ( .A1(n4855), .A2(n4832), .B1(n4457), .B2(n4854), .ZN(n2454)
         );
  AOI22_X1 U7323 ( .A1(n4857), .A2(n4832), .B1(n3937), .B2(n4856), .ZN(n2453)
         );
  AOI22_X1 U7324 ( .A1(n4859), .A2(n4832), .B1(n3938), .B2(n4858), .ZN(n2452)
         );
  AOI22_X1 U7325 ( .A1(n4861), .A2(n4832), .B1(n4458), .B2(n4860), .ZN(n2451)
         );
  AOI22_X1 U7326 ( .A1(n4863), .A2(n4832), .B1(n3939), .B2(n4862), .ZN(n2450)
         );
  AOI22_X1 U7327 ( .A1(n4865), .A2(n4832), .B1(n4459), .B2(n4864), .ZN(n2449)
         );
  AOI22_X1 U7328 ( .A1(n4867), .A2(n4832), .B1(n4226), .B2(n4866), .ZN(n2448)
         );
  AOI22_X1 U7329 ( .A1(n4869), .A2(n4832), .B1(n4227), .B2(n4868), .ZN(n2447)
         );
  AOI22_X1 U7330 ( .A1(n4871), .A2(n4832), .B1(n4460), .B2(n4870), .ZN(n2446)
         );
  AOI22_X1 U7331 ( .A1(n4873), .A2(n4832), .B1(n3940), .B2(n4872), .ZN(n2445)
         );
  AOI22_X1 U7332 ( .A1(n4875), .A2(n4832), .B1(n3941), .B2(n4874), .ZN(n2444)
         );
  AOI22_X1 U7333 ( .A1(n4877), .A2(n4832), .B1(n4461), .B2(n4876), .ZN(n2443)
         );
  AOI22_X1 U7334 ( .A1(n4879), .A2(n4832), .B1(n3942), .B2(n4878), .ZN(n2442)
         );
  AOI22_X1 U7335 ( .A1(n4881), .A2(n4832), .B1(n4462), .B2(n4880), .ZN(n2441)
         );
  AOI22_X1 U7336 ( .A1(n4883), .A2(n4832), .B1(n4228), .B2(n4882), .ZN(n2440)
         );
  AOI22_X1 U7337 ( .A1(n4885), .A2(n4832), .B1(n4229), .B2(n4884), .ZN(n2439)
         );
  AOI22_X1 U7338 ( .A1(n4887), .A2(n4832), .B1(n4463), .B2(n4886), .ZN(n2438)
         );
  AOI22_X1 U7339 ( .A1(n4889), .A2(n7275), .B1(n3943), .B2(n4888), .ZN(n2437)
         );
  AOI22_X1 U7340 ( .A1(n4891), .A2(n7275), .B1(n3944), .B2(n4890), .ZN(n2436)
         );
  AOI22_X1 U7341 ( .A1(n4893), .A2(n7275), .B1(n4464), .B2(n4892), .ZN(n2435)
         );
  AOI22_X1 U7342 ( .A1(n7978), .A2(n7275), .B1(n3945), .B2(n4894), .ZN(n2434)
         );
  AOI22_X1 U7343 ( .A1(n7979), .A2(n7275), .B1(n4465), .B2(n4896), .ZN(n2433)
         );
  AOI22_X1 U7344 ( .A1(n7980), .A2(n7275), .B1(n4230), .B2(n4898), .ZN(n2432)
         );
  AOI22_X1 U7345 ( .A1(n7981), .A2(n4832), .B1(n4231), .B2(n4900), .ZN(n2431)
         );
  AOI22_X1 U7346 ( .A1(n7982), .A2(n4832), .B1(n4466), .B2(n4902), .ZN(n2430)
         );
  AOI22_X1 U7347 ( .A1(n7983), .A2(n4832), .B1(n3946), .B2(n4904), .ZN(n2429)
         );
  AOI22_X1 U7348 ( .A1(n7984), .A2(n4832), .B1(n3947), .B2(n4906), .ZN(n2428)
         );
  AOI22_X1 U7349 ( .A1(n7985), .A2(n4832), .B1(n4467), .B2(n4908), .ZN(n2427)
         );
  NAND4_X1 U7350 ( .A1(n7279), .A2(n7278), .A3(n7277), .A4(n7276), .ZN(n7426)
         );
  INV_X1 U7351 ( .A(n7426), .ZN(n7621) );
  INV_X1 U7352 ( .A(n7521), .ZN(n7281) );
  OAI222_X1 U7353 ( .A1(n7427), .A2(n7621), .B1(n7282), .B2(n7281), .C1(n3772), 
        .C2(n7280), .ZN(n7738) );
  NAND2_X1 U7354 ( .A1(n7429), .A2(n7427), .ZN(n7388) );
  OAI21_X1 U7355 ( .B1(n7427), .B2(n7411), .A(n7388), .ZN(n7736) );
  OAI21_X1 U7356 ( .B1(alu_a_q[12]), .B2(n7872), .A(alu_b_q[12]), .ZN(n7297)
         );
  INV_X1 U7357 ( .A(n7297), .ZN(n7283) );
  AOI22_X1 U7358 ( .A1(n7356), .A2(n7410), .B1(n7342), .B2(n7283), .ZN(n7288)
         );
  NOR2_X1 U7359 ( .A1(n7878), .A2(n7389), .ZN(n7286) );
  OAI22_X1 U7360 ( .A1(n7284), .A2(n7383), .B1(n3777), .B2(n7867), .ZN(n7285)
         );
  AOI211_X1 U7361 ( .C1(n7874), .C2(n7413), .A(n7286), .B(n7285), .ZN(n7287)
         );
  OAI211_X1 U7362 ( .C1(n7430), .C2(n7736), .A(n7288), .B(n7287), .ZN(n7300)
         );
  NAND2_X1 U7363 ( .A1(n7892), .A2(n7290), .ZN(n7897) );
  AOI22_X1 U7364 ( .A1(n3352), .A2(n7302), .B1(n3353), .B2(n7303), .ZN(n7298)
         );
  NAND2_X1 U7365 ( .A1(n3777), .A2(n3806), .ZN(n7296) );
  NOR2_X1 U7366 ( .A1(n3777), .A2(alu_b_q[12]), .ZN(n7333) );
  NOR2_X1 U7367 ( .A1(alu_a_q[12]), .A2(n3806), .ZN(n7903) );
  OAI22_X1 U7368 ( .A1(n7303), .A2(n3842), .B1(n3764), .B2(n7302), .ZN(n7294)
         );
  OAI22_X1 U7369 ( .A1(n7333), .A2(n7903), .B1(n7835), .B2(n7294), .ZN(n7295)
         );
  OAI221_X1 U7370 ( .B1(n7298), .B2(n7297), .C1(n7298), .C2(n7296), .A(n7295), 
        .ZN(n7299) );
  AOI22_X1 U7371 ( .A1(n4847), .A2(n4833), .B1(n3948), .B2(n4846), .ZN(n2426)
         );
  AOI22_X1 U7372 ( .A1(n4849), .A2(n4833), .B1(n4468), .B2(n4848), .ZN(n2425)
         );
  AOI22_X1 U7373 ( .A1(n4851), .A2(n4833), .B1(n4232), .B2(n4850), .ZN(n2424)
         );
  AOI22_X1 U7374 ( .A1(n4853), .A2(n4833), .B1(n4233), .B2(n4852), .ZN(n2423)
         );
  AOI22_X1 U7375 ( .A1(n4855), .A2(n4833), .B1(n4469), .B2(n4854), .ZN(n2422)
         );
  AOI22_X1 U7376 ( .A1(n4857), .A2(n4833), .B1(n3949), .B2(n4856), .ZN(n2421)
         );
  AOI22_X1 U7377 ( .A1(n4859), .A2(n4833), .B1(n3950), .B2(n4858), .ZN(n2420)
         );
  AOI22_X1 U7378 ( .A1(n4861), .A2(n4833), .B1(n4470), .B2(n4860), .ZN(n2419)
         );
  AOI22_X1 U7379 ( .A1(n4863), .A2(n4833), .B1(n3951), .B2(n4862), .ZN(n2418)
         );
  AOI22_X1 U7380 ( .A1(n4865), .A2(n4833), .B1(n4471), .B2(n4864), .ZN(n2417)
         );
  AOI22_X1 U7381 ( .A1(n4867), .A2(n4833), .B1(n4234), .B2(n4866), .ZN(n2416)
         );
  AOI22_X1 U7382 ( .A1(n4869), .A2(n4833), .B1(n4235), .B2(n4868), .ZN(n2415)
         );
  AOI22_X1 U7383 ( .A1(n4871), .A2(n4833), .B1(n4472), .B2(n4870), .ZN(n2414)
         );
  AOI22_X1 U7384 ( .A1(n4873), .A2(n4833), .B1(n3952), .B2(n4872), .ZN(n2413)
         );
  AOI22_X1 U7385 ( .A1(n4875), .A2(n4833), .B1(n3953), .B2(n4874), .ZN(n2412)
         );
  AOI22_X1 U7386 ( .A1(n4877), .A2(n4833), .B1(n4473), .B2(n4876), .ZN(n2411)
         );
  AOI22_X1 U7387 ( .A1(n4879), .A2(n4833), .B1(n3954), .B2(n4878), .ZN(n2410)
         );
  AOI22_X1 U7388 ( .A1(n4881), .A2(n4833), .B1(n4474), .B2(n4880), .ZN(n2409)
         );
  AOI22_X1 U7389 ( .A1(n4883), .A2(n4833), .B1(n4236), .B2(n4882), .ZN(n2408)
         );
  AOI22_X1 U7390 ( .A1(n4885), .A2(n4833), .B1(n4237), .B2(n4884), .ZN(n2407)
         );
  AOI22_X1 U7391 ( .A1(n4887), .A2(n4833), .B1(n4475), .B2(n4886), .ZN(n2406)
         );
  AOI22_X1 U7392 ( .A1(n4889), .A2(n7301), .B1(n3955), .B2(n4888), .ZN(n2405)
         );
  AOI22_X1 U7393 ( .A1(n4891), .A2(n7301), .B1(n3956), .B2(n4890), .ZN(n2404)
         );
  AOI22_X1 U7394 ( .A1(n4893), .A2(n7301), .B1(n4476), .B2(n4892), .ZN(n2403)
         );
  AOI22_X1 U7395 ( .A1(n7978), .A2(n7301), .B1(n3957), .B2(n4894), .ZN(n2402)
         );
  AOI22_X1 U7396 ( .A1(n7979), .A2(n7301), .B1(n4477), .B2(n4896), .ZN(n2401)
         );
  AOI22_X1 U7397 ( .A1(n7980), .A2(n7301), .B1(n4238), .B2(n4898), .ZN(n2400)
         );
  AOI22_X1 U7398 ( .A1(n7981), .A2(n4833), .B1(n4239), .B2(n4900), .ZN(n2399)
         );
  AOI22_X1 U7399 ( .A1(n7982), .A2(n4833), .B1(n4478), .B2(n4902), .ZN(n2398)
         );
  AOI22_X1 U7400 ( .A1(n7983), .A2(n4833), .B1(n3958), .B2(n4904), .ZN(n2397)
         );
  AOI22_X1 U7401 ( .A1(n7984), .A2(n4833), .B1(n3959), .B2(n4906), .ZN(n2396)
         );
  AOI22_X1 U7402 ( .A1(n7985), .A2(n4833), .B1(n4479), .B2(n4908), .ZN(n2395)
         );
  NOR2_X1 U7403 ( .A1(alu_a_q[13]), .A2(alu_b_q[13]), .ZN(n7336) );
  NOR2_X1 U7404 ( .A1(n7333), .A2(n7335), .ZN(n7323) );
  INV_X1 U7405 ( .A(n7323), .ZN(n7305) );
  NOR2_X1 U7406 ( .A1(n3777), .A2(n3806), .ZN(n7304) );
  OAI22_X1 U7407 ( .A1(n3764), .A2(n7305), .B1(n3842), .B2(n7337), .ZN(n7331)
         );
  OAI22_X1 U7408 ( .A1(n7307), .A2(n7391), .B1(n7306), .B2(n7385), .ZN(n7318)
         );
  NAND4_X1 U7409 ( .A1(n7311), .A2(n7310), .A3(n7309), .A4(n7308), .ZN(n7654)
         );
  AOI22_X1 U7410 ( .A1(n7414), .A2(n7654), .B1(n7424), .B2(n7552), .ZN(n7312)
         );
  OAI21_X1 U7411 ( .B1(n7314), .B2(n7313), .A(n7312), .ZN(n7315) );
  AOI21_X1 U7412 ( .B1(n7418), .B2(n7446), .A(n7315), .ZN(n7773) );
  OAI21_X1 U7413 ( .B1(n7427), .B2(n7316), .A(n7388), .ZN(n7786) );
  OAI22_X1 U7414 ( .A1(n7773), .A2(n7399), .B1(n7430), .B2(n7786), .ZN(n7317)
         );
  AOI211_X1 U7415 ( .C1(alu_a_q[13]), .C2(n7802), .A(n7318), .B(n7317), .ZN(
        n7321) );
  NAND2_X1 U7416 ( .A1(n7885), .A2(n7319), .ZN(n7320) );
  OAI211_X1 U7417 ( .C1(n7322), .C2(n7383), .A(n7321), .B(n7320), .ZN(n7330)
         );
  OAI21_X1 U7418 ( .B1(n7323), .B2(n3764), .A(n7865), .ZN(n7324) );
  AOI21_X1 U7419 ( .B1(n3353), .B2(n7337), .A(n7324), .ZN(n7328) );
  NAND2_X1 U7420 ( .A1(alu_a_q[13]), .A2(n7735), .ZN(n7325) );
  OAI21_X1 U7421 ( .B1(n7331), .B2(n7325), .A(alu_b_q[13]), .ZN(n7327) );
  NOR2_X1 U7422 ( .A1(alu_a_q[13]), .A2(n7872), .ZN(n7326) );
  NAND2_X1 U7423 ( .A1(alu_a_q[13]), .A2(n3776), .ZN(n7902) );
  AOI222_X1 U7424 ( .A1(n7328), .A2(n7327), .B1(n7328), .B2(n7326), .C1(n7327), 
        .C2(n7902), .ZN(n7329) );
  AOI22_X1 U7425 ( .A1(n4847), .A2(n4834), .B1(n3960), .B2(n4846), .ZN(n2394)
         );
  AOI22_X1 U7426 ( .A1(n4849), .A2(n4834), .B1(n4480), .B2(n4848), .ZN(n2393)
         );
  AOI22_X1 U7427 ( .A1(n4851), .A2(n4834), .B1(n4240), .B2(n4850), .ZN(n2392)
         );
  AOI22_X1 U7428 ( .A1(n4853), .A2(n4834), .B1(n4241), .B2(n4852), .ZN(n2391)
         );
  AOI22_X1 U7429 ( .A1(n4855), .A2(n4834), .B1(n4481), .B2(n4854), .ZN(n2390)
         );
  AOI22_X1 U7430 ( .A1(n4857), .A2(n4834), .B1(n3961), .B2(n4856), .ZN(n2389)
         );
  AOI22_X1 U7431 ( .A1(n4859), .A2(n4834), .B1(n3962), .B2(n4858), .ZN(n2388)
         );
  AOI22_X1 U7432 ( .A1(n4861), .A2(n4834), .B1(n4482), .B2(n4860), .ZN(n2387)
         );
  AOI22_X1 U7433 ( .A1(n4863), .A2(n4834), .B1(n3963), .B2(n4862), .ZN(n2386)
         );
  AOI22_X1 U7434 ( .A1(n4865), .A2(n4834), .B1(n4483), .B2(n4864), .ZN(n2385)
         );
  AOI22_X1 U7435 ( .A1(n4867), .A2(n4834), .B1(n4242), .B2(n4866), .ZN(n2384)
         );
  AOI22_X1 U7436 ( .A1(n4869), .A2(n7332), .B1(n4243), .B2(n4868), .ZN(n2383)
         );
  AOI22_X1 U7437 ( .A1(n4871), .A2(n4834), .B1(n4484), .B2(n4870), .ZN(n2382)
         );
  AOI22_X1 U7438 ( .A1(n4873), .A2(n4834), .B1(n3964), .B2(n4872), .ZN(n2381)
         );
  AOI22_X1 U7439 ( .A1(n4875), .A2(n7332), .B1(n3965), .B2(n4874), .ZN(n2380)
         );
  AOI22_X1 U7440 ( .A1(n4877), .A2(n7332), .B1(n4485), .B2(n4876), .ZN(n2379)
         );
  AOI22_X1 U7441 ( .A1(n4879), .A2(n7332), .B1(n3966), .B2(n4878), .ZN(n2378)
         );
  AOI22_X1 U7442 ( .A1(n4881), .A2(n7332), .B1(n4486), .B2(n4880), .ZN(n2377)
         );
  AOI22_X1 U7443 ( .A1(n4883), .A2(n7332), .B1(n4244), .B2(n4882), .ZN(n2376)
         );
  AOI22_X1 U7444 ( .A1(n4885), .A2(n4834), .B1(n4245), .B2(n4884), .ZN(n2375)
         );
  AOI22_X1 U7445 ( .A1(n4887), .A2(n4834), .B1(n4487), .B2(n4886), .ZN(n2374)
         );
  AOI22_X1 U7446 ( .A1(n4889), .A2(n4834), .B1(n3967), .B2(n4888), .ZN(n2373)
         );
  AOI22_X1 U7447 ( .A1(n4891), .A2(n4834), .B1(n3968), .B2(n4890), .ZN(n2372)
         );
  AOI22_X1 U7448 ( .A1(n4893), .A2(n4834), .B1(n4488), .B2(n4892), .ZN(n2371)
         );
  AOI22_X1 U7449 ( .A1(n7978), .A2(n4834), .B1(n3969), .B2(n4894), .ZN(n2370)
         );
  AOI22_X1 U7450 ( .A1(n7979), .A2(n4834), .B1(n4489), .B2(n4896), .ZN(n2369)
         );
  AOI22_X1 U7451 ( .A1(n7980), .A2(n4834), .B1(n4246), .B2(n4898), .ZN(n2368)
         );
  AOI22_X1 U7452 ( .A1(n7981), .A2(n4834), .B1(n4247), .B2(n4900), .ZN(n2367)
         );
  AOI22_X1 U7453 ( .A1(n7982), .A2(n4834), .B1(n4490), .B2(n4902), .ZN(n2366)
         );
  AOI22_X1 U7454 ( .A1(n7983), .A2(n4834), .B1(n3970), .B2(n4904), .ZN(n2365)
         );
  AOI22_X1 U7455 ( .A1(n7984), .A2(n4834), .B1(n3971), .B2(n4906), .ZN(n2364)
         );
  AOI22_X1 U7456 ( .A1(n7985), .A2(n4834), .B1(n4491), .B2(n4908), .ZN(n2363)
         );
  INV_X1 U7457 ( .A(n7333), .ZN(n7334) );
  NAND2_X1 U7458 ( .A1(n7902), .A2(n7334), .ZN(n7895) );
  NOR2_X1 U7459 ( .A1(alu_a_q[14]), .A2(n3846), .ZN(n7901) );
  NAND2_X1 U7460 ( .A1(alu_a_q[14]), .A2(n3846), .ZN(n7407) );
  NOR2_X1 U7461 ( .A1(n7835), .A2(n7407), .ZN(n7338) );
  OAI222_X1 U7462 ( .A1(n7366), .A2(n3764), .B1(n7901), .B2(n7338), .C1(n3842), 
        .C2(n7368), .ZN(n7364) );
  NOR2_X1 U7463 ( .A1(alu_a_q[14]), .A2(alu_b_q[14]), .ZN(n7340) );
  AOI22_X1 U7464 ( .A1(n3352), .A2(n7366), .B1(n3353), .B2(n7368), .ZN(n7339)
         );
  OAI21_X1 U7465 ( .B1(n7340), .B2(n7369), .A(n7339), .ZN(n7363) );
  OAI21_X1 U7466 ( .B1(n7427), .B2(n7341), .A(n7388), .ZN(n7799) );
  AOI22_X1 U7467 ( .A1(n7624), .A2(n7901), .B1(n7369), .B2(n7342), .ZN(n7344)
         );
  NAND2_X1 U7468 ( .A1(alu_a_q[14]), .A2(n7802), .ZN(n7343) );
  OAI211_X1 U7469 ( .C1(n7799), .C2(n7430), .A(n7344), .B(n7343), .ZN(n7362)
         );
  INV_X1 U7470 ( .A(n7478), .ZN(n7350) );
  NAND4_X1 U7471 ( .A1(n7348), .A2(n7347), .A3(n7346), .A4(n7345), .ZN(n7679)
         );
  AOI22_X1 U7472 ( .A1(n7414), .A2(n7679), .B1(n7424), .B2(n7581), .ZN(n7349)
         );
  OAI21_X1 U7473 ( .B1(n7350), .B2(n7379), .A(n7349), .ZN(n7351) );
  AOI21_X1 U7474 ( .B1(n7417), .B2(n7479), .A(n7351), .ZN(n7812) );
  INV_X1 U7475 ( .A(n7352), .ZN(n7353) );
  AOI22_X1 U7476 ( .A1(n7356), .A2(n7355), .B1(n7354), .B2(n7353), .ZN(n7360)
         );
  AOI22_X1 U7477 ( .A1(n7885), .A2(n7358), .B1(n7874), .B2(n7357), .ZN(n7359)
         );
  OAI211_X1 U7478 ( .C1(n7812), .C2(n7399), .A(n7360), .B(n7359), .ZN(n7361)
         );
  AOI22_X1 U7479 ( .A1(n4847), .A2(n4835), .B1(n3972), .B2(n4846), .ZN(n2362)
         );
  AOI22_X1 U7480 ( .A1(n4849), .A2(n4835), .B1(n4492), .B2(n4848), .ZN(n2361)
         );
  AOI22_X1 U7481 ( .A1(n4851), .A2(n4835), .B1(n4248), .B2(n4850), .ZN(n2360)
         );
  AOI22_X1 U7482 ( .A1(n4853), .A2(n4835), .B1(n4249), .B2(n4852), .ZN(n2359)
         );
  AOI22_X1 U7483 ( .A1(n4855), .A2(n4835), .B1(n4493), .B2(n4854), .ZN(n2358)
         );
  AOI22_X1 U7484 ( .A1(n4857), .A2(n4835), .B1(n3973), .B2(n4856), .ZN(n2357)
         );
  AOI22_X1 U7485 ( .A1(n4859), .A2(n4835), .B1(n3974), .B2(n4858), .ZN(n2356)
         );
  AOI22_X1 U7486 ( .A1(n4861), .A2(n4835), .B1(n4494), .B2(n4860), .ZN(n2355)
         );
  AOI22_X1 U7487 ( .A1(n4863), .A2(n4835), .B1(n3975), .B2(n4862), .ZN(n2354)
         );
  AOI22_X1 U7488 ( .A1(n4865), .A2(n4835), .B1(n4495), .B2(n4864), .ZN(n2353)
         );
  AOI22_X1 U7489 ( .A1(n4867), .A2(n4835), .B1(n4250), .B2(n4866), .ZN(n2352)
         );
  AOI22_X1 U7490 ( .A1(n4869), .A2(n4835), .B1(n4251), .B2(n4868), .ZN(n2351)
         );
  AOI22_X1 U7491 ( .A1(n4871), .A2(n4835), .B1(n4496), .B2(n4870), .ZN(n2350)
         );
  AOI22_X1 U7492 ( .A1(n4873), .A2(n4835), .B1(n3976), .B2(n4872), .ZN(n2349)
         );
  AOI22_X1 U7493 ( .A1(n4875), .A2(n4835), .B1(n3977), .B2(n4874), .ZN(n2348)
         );
  AOI22_X1 U7494 ( .A1(n4877), .A2(n4835), .B1(n4497), .B2(n4876), .ZN(n2347)
         );
  AOI22_X1 U7495 ( .A1(n4879), .A2(n4835), .B1(n3978), .B2(n4878), .ZN(n2346)
         );
  AOI22_X1 U7496 ( .A1(n4881), .A2(n4835), .B1(n4498), .B2(n4880), .ZN(n2345)
         );
  AOI22_X1 U7497 ( .A1(n4883), .A2(n4835), .B1(n4252), .B2(n4882), .ZN(n2344)
         );
  AOI22_X1 U7498 ( .A1(n4885), .A2(n4835), .B1(n4253), .B2(n4884), .ZN(n2343)
         );
  AOI22_X1 U7499 ( .A1(n4887), .A2(n4835), .B1(n4499), .B2(n4886), .ZN(n2342)
         );
  AOI22_X1 U7500 ( .A1(n4889), .A2(n7365), .B1(n3979), .B2(n4888), .ZN(n2341)
         );
  AOI22_X1 U7501 ( .A1(n4891), .A2(n7365), .B1(n3980), .B2(n4890), .ZN(n2340)
         );
  AOI22_X1 U7502 ( .A1(n4893), .A2(n7365), .B1(n4500), .B2(n4892), .ZN(n2339)
         );
  AOI22_X1 U7503 ( .A1(n7978), .A2(n7365), .B1(n3981), .B2(n4894), .ZN(n2338)
         );
  AOI22_X1 U7504 ( .A1(n7979), .A2(n7365), .B1(n4501), .B2(n4896), .ZN(n2337)
         );
  AOI22_X1 U7505 ( .A1(n7980), .A2(n7365), .B1(n4254), .B2(n4898), .ZN(n2336)
         );
  AOI22_X1 U7506 ( .A1(n7981), .A2(n4835), .B1(n4255), .B2(n4900), .ZN(n2335)
         );
  AOI22_X1 U7507 ( .A1(n7982), .A2(n4835), .B1(n4502), .B2(n4902), .ZN(n2334)
         );
  AOI22_X1 U7508 ( .A1(n7983), .A2(n4835), .B1(n3982), .B2(n4904), .ZN(n2333)
         );
  AOI22_X1 U7509 ( .A1(n7984), .A2(n4835), .B1(n3983), .B2(n4906), .ZN(n2332)
         );
  AOI22_X1 U7510 ( .A1(n7985), .A2(n4835), .B1(n4503), .B2(n4908), .ZN(n2331)
         );
  INV_X1 U7511 ( .A(n7408), .ZN(n7367) );
  NAND2_X1 U7512 ( .A1(n7407), .A2(n7367), .ZN(n7370) );
  AOI22_X1 U7513 ( .A1(n3352), .A2(n7370), .B1(n3353), .B2(n7405), .ZN(n7372)
         );
  AOI211_X1 U7514 ( .C1(n7372), .C2(n7865), .A(alu_b_q[15]), .B(n3785), .ZN(
        n7403) );
  OAI22_X1 U7515 ( .A1(n3764), .A2(n7370), .B1(n3842), .B2(n7405), .ZN(n7395)
         );
  INV_X1 U7516 ( .A(n7395), .ZN(n7371) );
  NAND2_X1 U7517 ( .A1(alu_a_q[15]), .A2(alu_b_q[15]), .ZN(n7406) );
  AOI21_X1 U7518 ( .B1(n7735), .B2(n7371), .A(n7406), .ZN(n7402) );
  NAND2_X1 U7519 ( .A1(alu_b_q[15]), .A2(n3785), .ZN(n7904) );
  AOI21_X1 U7520 ( .B1(n7372), .B2(n7676), .A(n7904), .ZN(n7401) );
  INV_X1 U7521 ( .A(n7373), .ZN(n7377) );
  NAND4_X1 U7522 ( .A1(n7377), .A2(n7376), .A3(n7375), .A4(n7374), .ZN(n7702)
         );
  AOI22_X1 U7523 ( .A1(n7417), .A2(n7596), .B1(n7424), .B2(n7700), .ZN(n7378)
         );
  OAI21_X1 U7524 ( .B1(n7380), .B2(n7379), .A(n7378), .ZN(n7381) );
  AOI21_X1 U7525 ( .B1(n7414), .B2(n7702), .A(n7381), .ZN(n7852) );
  OAI22_X1 U7526 ( .A1(n7385), .A2(n7384), .B1(n7383), .B2(n7382), .ZN(n7386)
         );
  INV_X1 U7527 ( .A(n7386), .ZN(n7398) );
  NOR2_X1 U7528 ( .A1(alu_a_q[15]), .A2(alu_b_q[15]), .ZN(n7396) );
  NAND2_X1 U7529 ( .A1(n7388), .A2(n7387), .ZN(n7830) );
  OAI22_X1 U7530 ( .A1(n7390), .A2(n7389), .B1(n7430), .B2(n7830), .ZN(n7394)
         );
  OAI22_X1 U7531 ( .A1(n7392), .A2(n7391), .B1(n3785), .B2(n7867), .ZN(n7393)
         );
  AOI211_X1 U7532 ( .C1(n7396), .C2(n7395), .A(n7394), .B(n7393), .ZN(n7397)
         );
  OAI211_X1 U7533 ( .C1(n7852), .C2(n7399), .A(n7398), .B(n7397), .ZN(n7400)
         );
  AOI22_X1 U7534 ( .A1(n4847), .A2(n3368), .B1(n3984), .B2(n4846), .ZN(n2330)
         );
  AOI22_X1 U7535 ( .A1(n4849), .A2(n3368), .B1(n4504), .B2(n4848), .ZN(n2329)
         );
  AOI22_X1 U7536 ( .A1(n4851), .A2(n3368), .B1(n4256), .B2(n4850), .ZN(n2328)
         );
  AOI22_X1 U7537 ( .A1(n4853), .A2(n3368), .B1(n4257), .B2(n4852), .ZN(n2327)
         );
  AOI22_X1 U7538 ( .A1(n4855), .A2(n3368), .B1(n4505), .B2(n4854), .ZN(n2326)
         );
  AOI22_X1 U7539 ( .A1(n4857), .A2(n3368), .B1(n3985), .B2(n4856), .ZN(n2325)
         );
  AOI22_X1 U7540 ( .A1(n4859), .A2(n3368), .B1(n3986), .B2(n4858), .ZN(n2324)
         );
  AOI22_X1 U7541 ( .A1(n4861), .A2(n3368), .B1(n4506), .B2(n4860), .ZN(n2323)
         );
  AOI22_X1 U7542 ( .A1(n4863), .A2(n3368), .B1(n3987), .B2(n4862), .ZN(n2322)
         );
  AOI22_X1 U7543 ( .A1(n4865), .A2(n3368), .B1(n4507), .B2(n4864), .ZN(n2321)
         );
  AOI22_X1 U7544 ( .A1(n4867), .A2(n3368), .B1(n4258), .B2(n4866), .ZN(n2320)
         );
  AOI22_X1 U7545 ( .A1(n4869), .A2(n3368), .B1(n4259), .B2(n4868), .ZN(n2319)
         );
  AOI22_X1 U7546 ( .A1(n4871), .A2(n7404), .B1(n4508), .B2(n4870), .ZN(n2318)
         );
  AOI22_X1 U7547 ( .A1(n4873), .A2(n3368), .B1(n3988), .B2(n4872), .ZN(n2317)
         );
  AOI22_X1 U7548 ( .A1(n4875), .A2(n3368), .B1(n3989), .B2(n4874), .ZN(n2316)
         );
  AOI22_X1 U7549 ( .A1(n4877), .A2(n3368), .B1(n4509), .B2(n4876), .ZN(n2315)
         );
  AOI22_X1 U7550 ( .A1(n4879), .A2(n3368), .B1(n3990), .B2(n4878), .ZN(n2314)
         );
  AOI22_X1 U7551 ( .A1(n4881), .A2(n3368), .B1(n4510), .B2(n4880), .ZN(n2313)
         );
  AOI22_X1 U7552 ( .A1(n4883), .A2(n3368), .B1(n4260), .B2(n4882), .ZN(n2312)
         );
  AOI22_X1 U7553 ( .A1(n4885), .A2(n3368), .B1(n4261), .B2(n4884), .ZN(n2311)
         );
  AOI22_X1 U7554 ( .A1(n4887), .A2(n3368), .B1(n4511), .B2(n4886), .ZN(n2310)
         );
  AOI22_X1 U7555 ( .A1(n4889), .A2(n3368), .B1(n3991), .B2(n4888), .ZN(n2309)
         );
  AOI22_X1 U7556 ( .A1(n4891), .A2(n3368), .B1(n3992), .B2(n4890), .ZN(n2308)
         );
  AOI22_X1 U7557 ( .A1(n4893), .A2(n3368), .B1(n4512), .B2(n4892), .ZN(n2307)
         );
  AOI22_X1 U7558 ( .A1(n7978), .A2(n3368), .B1(n3993), .B2(n4894), .ZN(n2306)
         );
  AOI22_X1 U7559 ( .A1(n7979), .A2(n3368), .B1(n4513), .B2(n4896), .ZN(n2305)
         );
  AOI22_X1 U7560 ( .A1(n7980), .A2(n3368), .B1(n4262), .B2(n4898), .ZN(n2304)
         );
  AOI22_X1 U7561 ( .A1(n7981), .A2(n3368), .B1(n4263), .B2(n4900), .ZN(n2303)
         );
  AOI22_X1 U7562 ( .A1(n7982), .A2(n3368), .B1(n4514), .B2(n4902), .ZN(n2302)
         );
  AOI22_X1 U7563 ( .A1(n7983), .A2(n3368), .B1(n3994), .B2(n4904), .ZN(n2301)
         );
  AOI22_X1 U7564 ( .A1(n7984), .A2(n3368), .B1(n3995), .B2(n4906), .ZN(n2300)
         );
  AOI22_X1 U7565 ( .A1(n7985), .A2(n3368), .B1(n4515), .B2(n4908), .ZN(n2299)
         );
  OAI21_X1 U7566 ( .B1(alu_b_q[15]), .B2(n3785), .A(n7407), .ZN(n7905) );
  OAI22_X1 U7567 ( .A1(n7443), .A2(n3842), .B1(n3764), .B2(n7458), .ZN(n7409)
         );
  NOR2_X1 U7568 ( .A1(n7835), .A2(n7409), .ZN(n7436) );
  NAND2_X1 U7569 ( .A1(alu_a_q[16]), .A2(n3848), .ZN(n7907) );
  NAND2_X1 U7570 ( .A1(n3793), .A2(alu_b_q[16]), .ZN(n7457) );
  AOI22_X1 U7571 ( .A1(n7418), .A2(n7411), .B1(n7424), .B2(n7410), .ZN(n7416)
         );
  AOI22_X1 U7572 ( .A1(n7414), .A2(n7413), .B1(n7417), .B2(n7412), .ZN(n7415)
         );
  NAND2_X1 U7573 ( .A1(n7416), .A2(n7415), .ZN(n7946) );
  NAND2_X1 U7574 ( .A1(n7425), .A2(n7417), .ZN(n7709) );
  NAND2_X1 U7575 ( .A1(n7425), .A2(n7418), .ZN(n7620) );
  AOI22_X1 U7576 ( .A1(n7796), .A2(n7521), .B1(n7808), .B2(n7419), .ZN(n7433)
         );
  NAND4_X1 U7577 ( .A1(n7423), .A2(n7422), .A3(n7421), .A4(n7420), .ZN(n7619)
         );
  NAND2_X1 U7578 ( .A1(n7425), .A2(n7424), .ZN(n7708) );
  AOI22_X1 U7579 ( .A1(n7866), .A2(n7619), .B1(n7801), .B2(n7426), .ZN(n7432)
         );
  NOR2_X1 U7580 ( .A1(n7427), .A2(n7851), .ZN(n7701) );
  AOI22_X1 U7581 ( .A1(alu_a_q[16]), .A2(n7802), .B1(n7428), .B2(n7701), .ZN(
        n7431) );
  NAND4_X1 U7582 ( .A1(n7433), .A2(n7432), .A3(n7431), .A4(n7797), .ZN(n7434)
         );
  AOI21_X1 U7583 ( .B1(n7699), .B2(n7946), .A(n7434), .ZN(n7435) );
  OAI221_X1 U7584 ( .B1(n7436), .B2(n7907), .C1(n7436), .C2(n7457), .A(n7435), 
        .ZN(n7441) );
  AOI22_X1 U7585 ( .A1(n3352), .A2(n7458), .B1(n3353), .B2(n7443), .ZN(n7439)
         );
  OAI21_X1 U7586 ( .B1(alu_a_q[16]), .B2(n7872), .A(alu_b_q[16]), .ZN(n7438)
         );
  NAND2_X1 U7587 ( .A1(n3793), .A2(n3848), .ZN(n7437) );
  AOI222_X1 U7588 ( .A1(n7439), .A2(n7438), .B1(n7439), .B2(n7735), .C1(n7438), 
        .C2(n7437), .ZN(n7440) );
  AOI22_X1 U7589 ( .A1(n7954), .A2(n4836), .B1(n3996), .B2(n4846), .ZN(n2298)
         );
  AOI22_X1 U7590 ( .A1(n7955), .A2(n4836), .B1(n4516), .B2(n4848), .ZN(n2297)
         );
  AOI22_X1 U7591 ( .A1(n7956), .A2(n4836), .B1(n4264), .B2(n4850), .ZN(n2296)
         );
  AOI22_X1 U7592 ( .A1(n7957), .A2(n4836), .B1(n4265), .B2(n4852), .ZN(n2295)
         );
  AOI22_X1 U7593 ( .A1(n7958), .A2(n4836), .B1(n4517), .B2(n4854), .ZN(n2294)
         );
  AOI22_X1 U7594 ( .A1(n7959), .A2(n4836), .B1(n3997), .B2(n4856), .ZN(n2293)
         );
  AOI22_X1 U7595 ( .A1(n7960), .A2(n4836), .B1(n3998), .B2(n4858), .ZN(n2292)
         );
  AOI22_X1 U7596 ( .A1(n7961), .A2(n4836), .B1(n4518), .B2(n4860), .ZN(n2291)
         );
  AOI22_X1 U7597 ( .A1(n7962), .A2(n4836), .B1(n3999), .B2(n4862), .ZN(n2290)
         );
  AOI22_X1 U7598 ( .A1(n7963), .A2(n4836), .B1(n4519), .B2(n4864), .ZN(n2289)
         );
  AOI22_X1 U7599 ( .A1(n7964), .A2(n4836), .B1(n4266), .B2(n4866), .ZN(n2288)
         );
  AOI22_X1 U7600 ( .A1(n7965), .A2(n4836), .B1(n4267), .B2(n4868), .ZN(n2287)
         );
  AOI22_X1 U7601 ( .A1(n7966), .A2(n4836), .B1(n4520), .B2(n4870), .ZN(n2286)
         );
  AOI22_X1 U7602 ( .A1(n7967), .A2(n4836), .B1(n4000), .B2(n4872), .ZN(n2285)
         );
  AOI22_X1 U7603 ( .A1(n7968), .A2(n4836), .B1(n4001), .B2(n4874), .ZN(n2284)
         );
  AOI22_X1 U7604 ( .A1(n7969), .A2(n4836), .B1(n4521), .B2(n4876), .ZN(n2283)
         );
  AOI22_X1 U7605 ( .A1(n7970), .A2(n4836), .B1(n4002), .B2(n4878), .ZN(n2282)
         );
  AOI22_X1 U7606 ( .A1(n7971), .A2(n7442), .B1(n4522), .B2(n4880), .ZN(n2281)
         );
  AOI22_X1 U7607 ( .A1(n7972), .A2(n7442), .B1(n4268), .B2(n4882), .ZN(n2280)
         );
  AOI22_X1 U7608 ( .A1(n7973), .A2(n7442), .B1(n4269), .B2(n4884), .ZN(n2279)
         );
  AOI22_X1 U7609 ( .A1(n7974), .A2(n7442), .B1(n4523), .B2(n4886), .ZN(n2278)
         );
  AOI22_X1 U7610 ( .A1(n7975), .A2(n7442), .B1(n4003), .B2(n4888), .ZN(n2277)
         );
  AOI22_X1 U7611 ( .A1(n7976), .A2(n7442), .B1(n4004), .B2(n4890), .ZN(n2276)
         );
  AOI22_X1 U7612 ( .A1(n7977), .A2(n7442), .B1(n4524), .B2(n4892), .ZN(n2275)
         );
  AOI22_X1 U7613 ( .A1(n4895), .A2(n7442), .B1(n4005), .B2(n4894), .ZN(n2274)
         );
  AOI22_X1 U7614 ( .A1(n4897), .A2(n7442), .B1(n4525), .B2(n4896), .ZN(n2273)
         );
  AOI22_X1 U7615 ( .A1(n4899), .A2(n7442), .B1(n4270), .B2(n4898), .ZN(n2272)
         );
  AOI22_X1 U7616 ( .A1(n4901), .A2(n7442), .B1(n4271), .B2(n4900), .ZN(n2271)
         );
  AOI22_X1 U7617 ( .A1(n4903), .A2(n7442), .B1(n4526), .B2(n4902), .ZN(n2270)
         );
  AOI22_X1 U7618 ( .A1(n4905), .A2(n4836), .B1(n4006), .B2(n4904), .ZN(n2269)
         );
  AOI22_X1 U7619 ( .A1(n4907), .A2(n4836), .B1(n4007), .B2(n4906), .ZN(n2268)
         );
  AOI22_X1 U7620 ( .A1(n4909), .A2(n4836), .B1(n4527), .B2(n4908), .ZN(n2267)
         );
  NOR2_X1 U7621 ( .A1(n3794), .A2(alu_b_q[17]), .ZN(n7462) );
  INV_X1 U7622 ( .A(n7462), .ZN(n7910) );
  NOR2_X1 U7623 ( .A1(n3847), .A2(alu_a_q[17]), .ZN(n7891) );
  INV_X1 U7624 ( .A(n7891), .ZN(n7459) );
  NOR2_X1 U7625 ( .A1(n3793), .A2(n3848), .ZN(n7444) );
  AOI21_X1 U7626 ( .B1(n3353), .B2(n7472), .A(n7835), .ZN(n7445) );
  AOI21_X1 U7627 ( .B1(n7910), .B2(n7459), .A(n7445), .ZN(n7470) );
  AOI22_X1 U7628 ( .A1(alu_b_q[17]), .A2(n7872), .B1(n7801), .B2(n7654), .ZN(
        n7456) );
  AOI21_X1 U7629 ( .B1(n7796), .B2(n7552), .A(n7833), .ZN(n7455) );
  AOI22_X1 U7630 ( .A1(alu_a_q[17]), .A2(n7802), .B1(n7701), .B2(n7446), .ZN(
        n7454) );
  INV_X1 U7631 ( .A(n7447), .ZN(n7451) );
  NOR4_X1 U7632 ( .A1(n7451), .A2(n7450), .A3(n7449), .A4(n7448), .ZN(n7779)
         );
  INV_X1 U7633 ( .A(n7779), .ZN(n7648) );
  AOI22_X1 U7634 ( .A1(n7808), .A2(n7452), .B1(n7866), .B2(n7648), .ZN(n7453)
         );
  NAND4_X1 U7635 ( .A1(n7456), .A2(n7455), .A3(n7454), .A4(n7453), .ZN(n7469)
         );
  INV_X1 U7636 ( .A(n7457), .ZN(n7890) );
  NOR2_X1 U7637 ( .A1(n7462), .A2(n7891), .ZN(n7461) );
  OAI22_X1 U7638 ( .A1(n7462), .A2(n7483), .B1(n7461), .B2(n7460), .ZN(n7463)
         );
  OAI22_X1 U7639 ( .A1(n7464), .A2(n7831), .B1(n3764), .B2(n7463), .ZN(n7468)
         );
  NAND2_X1 U7640 ( .A1(alu_a_q[17]), .A2(alu_b_q[17]), .ZN(n7473) );
  OR2_X1 U7641 ( .A1(n3842), .A2(n7472), .ZN(n7466) );
  NAND2_X1 U7642 ( .A1(n3794), .A2(n3847), .ZN(n7465) );
  AOI222_X1 U7643 ( .A1(n7473), .A2(n7466), .B1(n7473), .B2(n7465), .C1(n7466), 
        .C2(n7788), .ZN(n7467) );
  AOI22_X1 U7644 ( .A1(n7954), .A2(n3369), .B1(n4008), .B2(n4846), .ZN(n2266)
         );
  AOI22_X1 U7645 ( .A1(n7955), .A2(n3369), .B1(n4528), .B2(n4848), .ZN(n2265)
         );
  AOI22_X1 U7646 ( .A1(n7956), .A2(n3369), .B1(n4272), .B2(n4850), .ZN(n2264)
         );
  AOI22_X1 U7647 ( .A1(n7957), .A2(n3369), .B1(n4273), .B2(n4852), .ZN(n2263)
         );
  AOI22_X1 U7648 ( .A1(n7958), .A2(n3369), .B1(n4529), .B2(n4854), .ZN(n2262)
         );
  AOI22_X1 U7649 ( .A1(n7959), .A2(n3369), .B1(n4009), .B2(n4856), .ZN(n2261)
         );
  AOI22_X1 U7650 ( .A1(n7960), .A2(n3369), .B1(n4010), .B2(n4858), .ZN(n2260)
         );
  AOI22_X1 U7651 ( .A1(n7961), .A2(n3369), .B1(n4530), .B2(n4860), .ZN(n2259)
         );
  AOI22_X1 U7652 ( .A1(n7962), .A2(n3369), .B1(n4011), .B2(n4862), .ZN(n2258)
         );
  AOI22_X1 U7653 ( .A1(n7963), .A2(n3369), .B1(n4531), .B2(n4864), .ZN(n2257)
         );
  AOI22_X1 U7654 ( .A1(n7964), .A2(n3369), .B1(n4274), .B2(n4866), .ZN(n2256)
         );
  AOI22_X1 U7655 ( .A1(n7965), .A2(n3369), .B1(n4275), .B2(n4868), .ZN(n2255)
         );
  AOI22_X1 U7656 ( .A1(n7966), .A2(n7471), .B1(n4532), .B2(n4870), .ZN(n2254)
         );
  AOI22_X1 U7657 ( .A1(n7967), .A2(n3369), .B1(n4012), .B2(n4872), .ZN(n2253)
         );
  AOI22_X1 U7658 ( .A1(n7968), .A2(n3369), .B1(n4013), .B2(n4874), .ZN(n2252)
         );
  AOI22_X1 U7659 ( .A1(n7969), .A2(n3369), .B1(n4533), .B2(n4876), .ZN(n2251)
         );
  AOI22_X1 U7660 ( .A1(n7970), .A2(n3369), .B1(n4014), .B2(n4878), .ZN(n2250)
         );
  AOI22_X1 U7661 ( .A1(n7971), .A2(n3369), .B1(n4534), .B2(n4880), .ZN(n2249)
         );
  AOI22_X1 U7662 ( .A1(n7972), .A2(n3369), .B1(n4276), .B2(n4882), .ZN(n2248)
         );
  AOI22_X1 U7663 ( .A1(n7973), .A2(n3369), .B1(n4277), .B2(n4884), .ZN(n2247)
         );
  AOI22_X1 U7664 ( .A1(n7974), .A2(n3369), .B1(n4535), .B2(n4886), .ZN(n2246)
         );
  AOI22_X1 U7665 ( .A1(n7975), .A2(n3369), .B1(n4015), .B2(n4888), .ZN(n2245)
         );
  AOI22_X1 U7666 ( .A1(n7976), .A2(n3369), .B1(n4016), .B2(n4890), .ZN(n2244)
         );
  AOI22_X1 U7667 ( .A1(n7977), .A2(n3369), .B1(n4536), .B2(n4892), .ZN(n2243)
         );
  AOI22_X1 U7668 ( .A1(n4895), .A2(n3369), .B1(n4017), .B2(n4894), .ZN(n2242)
         );
  AOI22_X1 U7669 ( .A1(n4897), .A2(n3369), .B1(n4537), .B2(n4896), .ZN(n2241)
         );
  AOI22_X1 U7670 ( .A1(n4899), .A2(n3369), .B1(n4278), .B2(n4898), .ZN(n2240)
         );
  AOI22_X1 U7671 ( .A1(n4901), .A2(n3369), .B1(n4279), .B2(n4900), .ZN(n2239)
         );
  AOI22_X1 U7672 ( .A1(n4903), .A2(n3369), .B1(n4538), .B2(n4902), .ZN(n2238)
         );
  AOI22_X1 U7673 ( .A1(n4905), .A2(n3369), .B1(n4018), .B2(n4904), .ZN(n2237)
         );
  AOI22_X1 U7674 ( .A1(n4907), .A2(n3369), .B1(n4019), .B2(n4906), .ZN(n2236)
         );
  AOI22_X1 U7675 ( .A1(n4909), .A2(n3369), .B1(n4539), .B2(n4908), .ZN(n2235)
         );
  NAND2_X1 U7676 ( .A1(n3786), .A2(n3838), .ZN(n7495) );
  OAI21_X1 U7677 ( .B1(n3838), .B2(n3786), .A(n7495), .ZN(n7484) );
  AOI221_X1 U7678 ( .B1(n7496), .B2(n7865), .C1(n3842), .C2(n7865), .A(n7484), 
        .ZN(n7493) );
  NAND4_X1 U7679 ( .A1(n7477), .A2(n7476), .A3(n7475), .A4(n7474), .ZN(n7807)
         );
  AOI22_X1 U7680 ( .A1(n7701), .A2(n7478), .B1(n7866), .B2(n7807), .ZN(n7482)
         );
  AOI22_X1 U7681 ( .A1(alu_a_q[18]), .A2(n7802), .B1(n7801), .B2(n7679), .ZN(
        n7481) );
  AOI22_X1 U7682 ( .A1(n7796), .A2(n7581), .B1(n7808), .B2(n7479), .ZN(n7480)
         );
  NAND4_X1 U7683 ( .A1(n7482), .A2(n7481), .A3(n7480), .A4(n7797), .ZN(n7492)
         );
  XNOR2_X1 U7684 ( .A(n7509), .B(n7484), .ZN(n7485) );
  OAI22_X1 U7685 ( .A1(n7486), .A2(n7831), .B1(n3764), .B2(n7485), .ZN(n7491)
         );
  NAND2_X1 U7686 ( .A1(n3353), .A2(n7496), .ZN(n7488) );
  AOI22_X1 U7687 ( .A1(n3786), .A2(n7734), .B1(n7488), .B2(n7735), .ZN(n7487)
         );
  INV_X1 U7688 ( .A(n7487), .ZN(n7489) );
  OAI22_X1 U7689 ( .A1(n3838), .A2(n7489), .B1(n7495), .B2(n7488), .ZN(n7490)
         );
  AOI22_X1 U7690 ( .A1(n7954), .A2(n3367), .B1(n4020), .B2(n4846), .ZN(n2234)
         );
  AOI22_X1 U7691 ( .A1(n7955), .A2(n3367), .B1(n4540), .B2(n4848), .ZN(n2233)
         );
  AOI22_X1 U7692 ( .A1(n7956), .A2(n3367), .B1(n4280), .B2(n4850), .ZN(n2232)
         );
  AOI22_X1 U7693 ( .A1(n7957), .A2(n3367), .B1(n4281), .B2(n4852), .ZN(n2231)
         );
  AOI22_X1 U7694 ( .A1(n7958), .A2(n3367), .B1(n4541), .B2(n4854), .ZN(n2230)
         );
  AOI22_X1 U7695 ( .A1(n7959), .A2(n3367), .B1(n4021), .B2(n4856), .ZN(n2229)
         );
  AOI22_X1 U7696 ( .A1(n7960), .A2(n3367), .B1(n4022), .B2(n4858), .ZN(n2228)
         );
  AOI22_X1 U7697 ( .A1(n7961), .A2(n3367), .B1(n4542), .B2(n4860), .ZN(n2227)
         );
  AOI22_X1 U7698 ( .A1(n7962), .A2(n3367), .B1(n4023), .B2(n4862), .ZN(n2226)
         );
  AOI22_X1 U7699 ( .A1(n7963), .A2(n3367), .B1(n4543), .B2(n4864), .ZN(n2225)
         );
  AOI22_X1 U7700 ( .A1(n7964), .A2(n3367), .B1(n4282), .B2(n4866), .ZN(n2224)
         );
  AOI22_X1 U7701 ( .A1(n7965), .A2(n3367), .B1(n4283), .B2(n4868), .ZN(n2223)
         );
  AOI22_X1 U7702 ( .A1(n7966), .A2(n7494), .B1(n4544), .B2(n4870), .ZN(n2222)
         );
  AOI22_X1 U7703 ( .A1(n7967), .A2(n3367), .B1(n4024), .B2(n4872), .ZN(n2221)
         );
  AOI22_X1 U7704 ( .A1(n7968), .A2(n3367), .B1(n4025), .B2(n4874), .ZN(n2220)
         );
  AOI22_X1 U7705 ( .A1(n7969), .A2(n3367), .B1(n4545), .B2(n4876), .ZN(n2219)
         );
  AOI22_X1 U7706 ( .A1(n7970), .A2(n3367), .B1(n4026), .B2(n4878), .ZN(n2218)
         );
  AOI22_X1 U7707 ( .A1(n7971), .A2(n3367), .B1(n4546), .B2(n4880), .ZN(n2217)
         );
  AOI22_X1 U7708 ( .A1(n7972), .A2(n3367), .B1(n4284), .B2(n4882), .ZN(n2216)
         );
  AOI22_X1 U7709 ( .A1(n7973), .A2(n3367), .B1(n4285), .B2(n4884), .ZN(n2215)
         );
  AOI22_X1 U7710 ( .A1(n7974), .A2(n3367), .B1(n4547), .B2(n4886), .ZN(n2214)
         );
  AOI22_X1 U7711 ( .A1(n7975), .A2(n3367), .B1(n4027), .B2(n4888), .ZN(n2213)
         );
  AOI22_X1 U7712 ( .A1(n7976), .A2(n3367), .B1(n4028), .B2(n4890), .ZN(n2212)
         );
  AOI22_X1 U7713 ( .A1(n7977), .A2(n3367), .B1(n4548), .B2(n4892), .ZN(n2211)
         );
  AOI22_X1 U7714 ( .A1(n4895), .A2(n3367), .B1(n4029), .B2(n4894), .ZN(n2210)
         );
  AOI22_X1 U7715 ( .A1(n4897), .A2(n3367), .B1(n4549), .B2(n4896), .ZN(n2209)
         );
  AOI22_X1 U7716 ( .A1(n4899), .A2(n3367), .B1(n4286), .B2(n4898), .ZN(n2208)
         );
  AOI22_X1 U7717 ( .A1(n4901), .A2(n3367), .B1(n4287), .B2(n4900), .ZN(n2207)
         );
  AOI22_X1 U7718 ( .A1(n4903), .A2(n3367), .B1(n4550), .B2(n4902), .ZN(n2206)
         );
  AOI22_X1 U7719 ( .A1(n4905), .A2(n3367), .B1(n4030), .B2(n4904), .ZN(n2205)
         );
  AOI22_X1 U7720 ( .A1(n4907), .A2(n3367), .B1(n4031), .B2(n4906), .ZN(n2204)
         );
  AOI22_X1 U7721 ( .A1(n4909), .A2(n3367), .B1(n4551), .B2(n4908), .ZN(n2203)
         );
  NAND2_X1 U7722 ( .A1(alu_a_q[19]), .A2(n3850), .ZN(n7914) );
  NAND2_X1 U7723 ( .A1(alu_b_q[19]), .A2(n3787), .ZN(n7530) );
  OAI22_X1 U7724 ( .A1(n7735), .A2(n3787), .B1(n7532), .B2(n3842), .ZN(n7518)
         );
  NAND2_X1 U7725 ( .A1(n3353), .A2(n7532), .ZN(n7497) );
  AOI21_X1 U7726 ( .B1(n7865), .B2(n7497), .A(n7914), .ZN(n7517) );
  AOI21_X1 U7727 ( .B1(n3353), .B2(n7532), .A(n7624), .ZN(n7515) );
  AOI22_X1 U7728 ( .A1(n7498), .A2(n7701), .B1(n7702), .B2(n7801), .ZN(n7499)
         );
  INV_X1 U7729 ( .A(n7499), .ZN(n7508) );
  OAI22_X1 U7730 ( .A1(n7500), .A2(n7620), .B1(n3787), .B2(n7867), .ZN(n7507)
         );
  NOR4_X1 U7731 ( .A1(n7504), .A2(n7503), .A3(n7502), .A4(n7501), .ZN(n7842)
         );
  OAI22_X1 U7732 ( .A1(n7842), .A2(n7707), .B1(n7505), .B2(n7709), .ZN(n7506)
         );
  NOR4_X1 U7733 ( .A1(n7833), .A2(n7508), .A3(n7507), .A4(n7506), .ZN(n7514)
         );
  AOI21_X1 U7734 ( .B1(alu_b_q[18]), .B2(n3786), .A(n7531), .ZN(n7510) );
  XOR2_X1 U7735 ( .A(n7510), .B(n7519), .Z(n7512) );
  AOI22_X1 U7736 ( .A1(n3352), .A2(n7512), .B1(n7699), .B2(n7511), .ZN(n7513)
         );
  OAI211_X1 U7737 ( .C1(n7515), .C2(n7530), .A(n7514), .B(n7513), .ZN(n7516)
         );
  AOI22_X1 U7738 ( .A1(n7954), .A2(n4837), .B1(n4032), .B2(n4846), .ZN(n2202)
         );
  AOI22_X1 U7739 ( .A1(n7955), .A2(n4837), .B1(n4552), .B2(n4848), .ZN(n2201)
         );
  AOI22_X1 U7740 ( .A1(n7956), .A2(n4837), .B1(n4288), .B2(n4850), .ZN(n2200)
         );
  AOI22_X1 U7741 ( .A1(n7957), .A2(n4837), .B1(n4289), .B2(n4852), .ZN(n2199)
         );
  AOI22_X1 U7742 ( .A1(n7958), .A2(n4837), .B1(n4553), .B2(n4854), .ZN(n2198)
         );
  AOI22_X1 U7743 ( .A1(n7959), .A2(n4837), .B1(n4033), .B2(n4856), .ZN(n2197)
         );
  AOI22_X1 U7744 ( .A1(n7960), .A2(n4837), .B1(n4034), .B2(n4858), .ZN(n2196)
         );
  AOI22_X1 U7745 ( .A1(n7961), .A2(n4837), .B1(n4554), .B2(n4860), .ZN(n2195)
         );
  AOI22_X1 U7746 ( .A1(n7962), .A2(n4837), .B1(n4035), .B2(n4862), .ZN(n2194)
         );
  AOI22_X1 U7747 ( .A1(n7963), .A2(n4837), .B1(n4555), .B2(n4864), .ZN(n2193)
         );
  AOI22_X1 U7748 ( .A1(n7964), .A2(n4837), .B1(n4290), .B2(n4866), .ZN(n2192)
         );
  AOI22_X1 U7749 ( .A1(n7965), .A2(n4837), .B1(n4291), .B2(n4868), .ZN(n2191)
         );
  AOI22_X1 U7750 ( .A1(n7966), .A2(n4837), .B1(n4556), .B2(n4870), .ZN(n2190)
         );
  AOI22_X1 U7751 ( .A1(n7967), .A2(n4837), .B1(n4036), .B2(n4872), .ZN(n2189)
         );
  AOI22_X1 U7752 ( .A1(n7968), .A2(n4837), .B1(n4037), .B2(n4874), .ZN(n2188)
         );
  AOI22_X1 U7753 ( .A1(n7969), .A2(n4837), .B1(n4557), .B2(n4876), .ZN(n2187)
         );
  AOI22_X1 U7754 ( .A1(n7970), .A2(n4837), .B1(n4038), .B2(n4878), .ZN(n2186)
         );
  AOI22_X1 U7755 ( .A1(n7971), .A2(n4837), .B1(n4558), .B2(n4880), .ZN(n2185)
         );
  AOI22_X1 U7756 ( .A1(n7972), .A2(n4837), .B1(n4292), .B2(n4882), .ZN(n2184)
         );
  AOI22_X1 U7757 ( .A1(n7973), .A2(n4837), .B1(n4293), .B2(n4884), .ZN(n2183)
         );
  AOI22_X1 U7758 ( .A1(n7974), .A2(n4837), .B1(n4559), .B2(n4886), .ZN(n2182)
         );
  AOI22_X1 U7759 ( .A1(n7975), .A2(n7520), .B1(n4039), .B2(n4888), .ZN(n2181)
         );
  AOI22_X1 U7760 ( .A1(n7976), .A2(n7520), .B1(n4040), .B2(n4890), .ZN(n2180)
         );
  AOI22_X1 U7761 ( .A1(n7977), .A2(n7520), .B1(n4560), .B2(n4892), .ZN(n2179)
         );
  AOI22_X1 U7762 ( .A1(n4895), .A2(n7520), .B1(n4041), .B2(n4894), .ZN(n2178)
         );
  AOI22_X1 U7763 ( .A1(n4897), .A2(n7520), .B1(n4561), .B2(n4896), .ZN(n2177)
         );
  AOI22_X1 U7764 ( .A1(n4899), .A2(n7520), .B1(n4294), .B2(n4898), .ZN(n2176)
         );
  AOI22_X1 U7765 ( .A1(n4901), .A2(n4837), .B1(n4295), .B2(n4900), .ZN(n2175)
         );
  AOI22_X1 U7766 ( .A1(n4903), .A2(n4837), .B1(n4562), .B2(n4902), .ZN(n2174)
         );
  AOI22_X1 U7767 ( .A1(n4905), .A2(n4837), .B1(n4042), .B2(n4904), .ZN(n2173)
         );
  AOI22_X1 U7768 ( .A1(n4907), .A2(n4837), .B1(n4043), .B2(n4906), .ZN(n2172)
         );
  AOI22_X1 U7769 ( .A1(n4909), .A2(n4837), .B1(n4563), .B2(n4908), .ZN(n2171)
         );
  AOI22_X1 U7770 ( .A1(n7808), .A2(n7521), .B1(n7801), .B2(n7619), .ZN(n7528)
         );
  OAI22_X1 U7771 ( .A1(n7750), .A2(n7707), .B1(n7621), .B2(n7709), .ZN(n7526)
         );
  AOI211_X1 U7772 ( .C1(alu_a_q[20]), .C2(n7802), .A(n7833), .B(n7526), .ZN(
        n7527) );
  OAI211_X1 U7773 ( .C1(n7529), .C2(n7831), .A(n7528), .B(n7527), .ZN(n7543)
         );
  OAI21_X1 U7774 ( .B1(alu_a_q[18]), .B2(n3838), .A(n7530), .ZN(n7917) );
  AOI222_X1 U7775 ( .A1(n7532), .A2(n3850), .B1(n7532), .B2(n3787), .C1(n3850), 
        .C2(n3787), .ZN(n7557) );
  AOI22_X1 U7776 ( .A1(n3352), .A2(n7555), .B1(n3353), .B2(n7557), .ZN(n7541)
         );
  NAND2_X1 U7777 ( .A1(n3791), .A2(n3849), .ZN(n7556) );
  AND2_X1 U7778 ( .A1(alu_a_q[20]), .A2(n7541), .ZN(n7533) );
  AOI21_X1 U7779 ( .B1(n7533), .B2(n7735), .A(n3849), .ZN(n7539) );
  AOI21_X1 U7780 ( .B1(n3352), .B2(n7534), .A(n7835), .ZN(n7535) );
  OAI21_X1 U7781 ( .B1(n7557), .B2(n3842), .A(n7535), .ZN(n7538) );
  NAND2_X1 U7782 ( .A1(n3791), .A2(n7734), .ZN(n7537) );
  NAND2_X1 U7783 ( .A1(n3849), .A2(alu_a_q[20]), .ZN(n7915) );
  INV_X1 U7784 ( .A(n7915), .ZN(n7536) );
  AOI222_X1 U7785 ( .A1(n7539), .A2(n7538), .B1(n7539), .B2(n7537), .C1(n7538), 
        .C2(n7536), .ZN(n7540) );
  OAI21_X1 U7786 ( .B1(n7541), .B2(n7556), .A(n7540), .ZN(n7542) );
  AOI22_X1 U7787 ( .A1(n7954), .A2(n4838), .B1(n4044), .B2(n4846), .ZN(n2170)
         );
  AOI22_X1 U7788 ( .A1(n7955), .A2(n4838), .B1(n4564), .B2(n4848), .ZN(n2169)
         );
  AOI22_X1 U7789 ( .A1(n7956), .A2(n4838), .B1(n4296), .B2(n4850), .ZN(n2168)
         );
  AOI22_X1 U7790 ( .A1(n7957), .A2(n4838), .B1(n4297), .B2(n4852), .ZN(n2167)
         );
  AOI22_X1 U7791 ( .A1(n7958), .A2(n4838), .B1(n4565), .B2(n4854), .ZN(n2166)
         );
  AOI22_X1 U7792 ( .A1(n7959), .A2(n4838), .B1(n4045), .B2(n4856), .ZN(n2165)
         );
  AOI22_X1 U7793 ( .A1(n7960), .A2(n4838), .B1(n4046), .B2(n4858), .ZN(n2164)
         );
  AOI22_X1 U7794 ( .A1(n7961), .A2(n4838), .B1(n4566), .B2(n4860), .ZN(n2163)
         );
  AOI22_X1 U7795 ( .A1(n7962), .A2(n4838), .B1(n4047), .B2(n4862), .ZN(n2162)
         );
  AOI22_X1 U7796 ( .A1(n7963), .A2(n4838), .B1(n4567), .B2(n4864), .ZN(n2161)
         );
  AOI22_X1 U7797 ( .A1(n7964), .A2(n4838), .B1(n4298), .B2(n4866), .ZN(n2160)
         );
  AOI22_X1 U7798 ( .A1(n7965), .A2(n4838), .B1(n4299), .B2(n4868), .ZN(n2159)
         );
  AOI22_X1 U7799 ( .A1(n7966), .A2(n4838), .B1(n4568), .B2(n4870), .ZN(n2158)
         );
  AOI22_X1 U7800 ( .A1(n7967), .A2(n4838), .B1(n4048), .B2(n4872), .ZN(n2157)
         );
  AOI22_X1 U7801 ( .A1(n7968), .A2(n4838), .B1(n4049), .B2(n4874), .ZN(n2156)
         );
  AOI22_X1 U7802 ( .A1(n7969), .A2(n4838), .B1(n4569), .B2(n4876), .ZN(n2155)
         );
  AOI22_X1 U7803 ( .A1(n7970), .A2(n4838), .B1(n4050), .B2(n4878), .ZN(n2154)
         );
  AOI22_X1 U7804 ( .A1(n7971), .A2(n4838), .B1(n4570), .B2(n4880), .ZN(n2153)
         );
  AOI22_X1 U7805 ( .A1(n7972), .A2(n4838), .B1(n4300), .B2(n4882), .ZN(n2152)
         );
  AOI22_X1 U7806 ( .A1(n7973), .A2(n4838), .B1(n4301), .B2(n4884), .ZN(n2151)
         );
  AOI22_X1 U7807 ( .A1(n7974), .A2(n4838), .B1(n4571), .B2(n4886), .ZN(n2150)
         );
  AOI22_X1 U7808 ( .A1(n7975), .A2(n7545), .B1(n4051), .B2(n4888), .ZN(n2149)
         );
  AOI22_X1 U7809 ( .A1(n7976), .A2(n7545), .B1(n4052), .B2(n4890), .ZN(n2148)
         );
  AOI22_X1 U7810 ( .A1(n7977), .A2(n7545), .B1(n4572), .B2(n4892), .ZN(n2147)
         );
  AOI22_X1 U7811 ( .A1(n4895), .A2(n7545), .B1(n4053), .B2(n4894), .ZN(n2146)
         );
  AOI22_X1 U7812 ( .A1(n4897), .A2(n7545), .B1(n4573), .B2(n4896), .ZN(n2145)
         );
  AOI22_X1 U7813 ( .A1(n4899), .A2(n7545), .B1(n4302), .B2(n4898), .ZN(n2144)
         );
  AOI22_X1 U7814 ( .A1(n4901), .A2(n4838), .B1(n4303), .B2(n4900), .ZN(n2143)
         );
  AOI22_X1 U7815 ( .A1(n4903), .A2(n4838), .B1(n4574), .B2(n4902), .ZN(n2142)
         );
  AOI22_X1 U7816 ( .A1(n4905), .A2(n4838), .B1(n4054), .B2(n4904), .ZN(n2141)
         );
  AOI22_X1 U7817 ( .A1(n4907), .A2(n4838), .B1(n4055), .B2(n4906), .ZN(n2140)
         );
  AOI22_X1 U7818 ( .A1(n4909), .A2(n4838), .B1(n4575), .B2(n4908), .ZN(n2139)
         );
  AOI22_X1 U7819 ( .A1(alu_b_q[21]), .A2(n7872), .B1(n7801), .B2(n7648), .ZN(
        n7546) );
  OAI211_X1 U7820 ( .C1(n7547), .C2(n7851), .A(n7546), .B(n7797), .ZN(n7566)
         );
  NOR4_X1 U7821 ( .A1(n7551), .A2(n7550), .A3(n7549), .A4(n7548), .ZN(n7781)
         );
  OAI22_X1 U7822 ( .A1(n7781), .A2(n7707), .B1(n3766), .B2(n7867), .ZN(n7565)
         );
  AOI22_X1 U7823 ( .A1(n7796), .A2(n7654), .B1(n7808), .B2(n7552), .ZN(n7553)
         );
  OAI21_X1 U7824 ( .B1(n7554), .B2(n7831), .A(n7553), .ZN(n7564) );
  OAI221_X1 U7825 ( .B1(n7557), .B2(alu_b_q[20]), .C1(n7557), .C2(alu_a_q[20]), 
        .A(n7556), .ZN(n7574) );
  OAI222_X1 U7826 ( .A1(n7576), .A2(n3764), .B1(n3842), .B2(n7574), .C1(n3839), 
        .C2(n7788), .ZN(n7558) );
  INV_X1 U7827 ( .A(n7558), .ZN(n7562) );
  NAND2_X1 U7828 ( .A1(alu_a_q[21]), .A2(alu_b_q[21]), .ZN(n7575) );
  OAI21_X1 U7829 ( .B1(alu_a_q[21]), .B2(alu_b_q[21]), .A(n7575), .ZN(n7561)
         );
  AOI22_X1 U7830 ( .A1(n3352), .A2(n7576), .B1(n3353), .B2(n7574), .ZN(n7560)
         );
  NOR2_X1 U7831 ( .A1(n7561), .A2(n7835), .ZN(n7559) );
  AOI22_X1 U7832 ( .A1(n7562), .A2(n7561), .B1(n7560), .B2(n7559), .ZN(n7563)
         );
  AOI22_X1 U7833 ( .A1(n4847), .A2(n3366), .B1(n4056), .B2(n4846), .ZN(n2138)
         );
  AOI22_X1 U7834 ( .A1(n4849), .A2(n3366), .B1(n4576), .B2(n4848), .ZN(n2137)
         );
  AOI22_X1 U7835 ( .A1(n4851), .A2(n3366), .B1(n4304), .B2(n4850), .ZN(n2136)
         );
  AOI22_X1 U7836 ( .A1(n4853), .A2(n3366), .B1(n4305), .B2(n4852), .ZN(n2135)
         );
  AOI22_X1 U7837 ( .A1(n4855), .A2(n3366), .B1(n4577), .B2(n4854), .ZN(n2134)
         );
  AOI22_X1 U7838 ( .A1(n4857), .A2(n3366), .B1(n4057), .B2(n4856), .ZN(n2133)
         );
  AOI22_X1 U7839 ( .A1(n4859), .A2(n3366), .B1(n4058), .B2(n4858), .ZN(n2132)
         );
  AOI22_X1 U7840 ( .A1(n4861), .A2(n3366), .B1(n4578), .B2(n4860), .ZN(n2131)
         );
  AOI22_X1 U7841 ( .A1(n4863), .A2(n3366), .B1(n4059), .B2(n4862), .ZN(n2130)
         );
  AOI22_X1 U7842 ( .A1(n4865), .A2(n3366), .B1(n4579), .B2(n4864), .ZN(n2129)
         );
  AOI22_X1 U7843 ( .A1(n4867), .A2(n3366), .B1(n4306), .B2(n4866), .ZN(n2128)
         );
  AOI22_X1 U7844 ( .A1(n4869), .A2(n3366), .B1(n4307), .B2(n4868), .ZN(n2127)
         );
  AOI22_X1 U7845 ( .A1(n4871), .A2(n7567), .B1(n4580), .B2(n4870), .ZN(n2126)
         );
  AOI22_X1 U7846 ( .A1(n4873), .A2(n3366), .B1(n4060), .B2(n4872), .ZN(n2125)
         );
  AOI22_X1 U7847 ( .A1(n4875), .A2(n3366), .B1(n4061), .B2(n4874), .ZN(n2124)
         );
  AOI22_X1 U7848 ( .A1(n4877), .A2(n3366), .B1(n4581), .B2(n4876), .ZN(n2123)
         );
  AOI22_X1 U7849 ( .A1(n4879), .A2(n3366), .B1(n4062), .B2(n4878), .ZN(n2122)
         );
  AOI22_X1 U7850 ( .A1(n4881), .A2(n3366), .B1(n4582), .B2(n4880), .ZN(n2121)
         );
  AOI22_X1 U7851 ( .A1(n4883), .A2(n3366), .B1(n4308), .B2(n4882), .ZN(n2120)
         );
  AOI22_X1 U7852 ( .A1(n4885), .A2(n3366), .B1(n4309), .B2(n4884), .ZN(n2119)
         );
  AOI22_X1 U7853 ( .A1(n4887), .A2(n3366), .B1(n4583), .B2(n4886), .ZN(n2118)
         );
  AOI22_X1 U7854 ( .A1(n4889), .A2(n3366), .B1(n4063), .B2(n4888), .ZN(n2117)
         );
  AOI22_X1 U7855 ( .A1(n4891), .A2(n3366), .B1(n4064), .B2(n4890), .ZN(n2116)
         );
  AOI22_X1 U7856 ( .A1(n4893), .A2(n3366), .B1(n4584), .B2(n4892), .ZN(n2115)
         );
  AOI22_X1 U7857 ( .A1(n4895), .A2(n3366), .B1(n4065), .B2(n4894), .ZN(n2114)
         );
  AOI22_X1 U7858 ( .A1(n4897), .A2(n3366), .B1(n4585), .B2(n4896), .ZN(n2113)
         );
  AOI22_X1 U7859 ( .A1(n4899), .A2(n3366), .B1(n4310), .B2(n4898), .ZN(n2112)
         );
  AOI22_X1 U7860 ( .A1(n4901), .A2(n3366), .B1(n4311), .B2(n4900), .ZN(n2111)
         );
  AOI22_X1 U7861 ( .A1(n4903), .A2(n3366), .B1(n4586), .B2(n4902), .ZN(n2110)
         );
  AOI22_X1 U7862 ( .A1(n4905), .A2(n3366), .B1(n4066), .B2(n4904), .ZN(n2109)
         );
  AOI22_X1 U7863 ( .A1(n4907), .A2(n3366), .B1(n4067), .B2(n4906), .ZN(n2108)
         );
  AOI22_X1 U7864 ( .A1(n4909), .A2(n3366), .B1(n4587), .B2(n4908), .ZN(n2107)
         );
  NAND4_X1 U7865 ( .A1(n7571), .A2(n7570), .A3(n7569), .A4(n7568), .ZN(n7795)
         );
  AOI22_X1 U7866 ( .A1(alu_b_q[22]), .A2(n7872), .B1(n7866), .B2(n7795), .ZN(
        n7572) );
  OAI211_X1 U7867 ( .C1(n7573), .C2(n7851), .A(n7572), .B(n7797), .ZN(n7587)
         );
  NOR2_X1 U7868 ( .A1(n3795), .A2(n3845), .ZN(n7591) );
  NAND2_X1 U7869 ( .A1(n7591), .A2(n7788), .ZN(n7577) );
  NOR2_X1 U7870 ( .A1(alu_a_q[22]), .A2(alu_b_q[22]), .ZN(n7580) );
  INV_X1 U7871 ( .A(n7580), .ZN(n7592) );
  NOR2_X1 U7872 ( .A1(n3766), .A2(alu_b_q[21]), .ZN(n7921) );
  OAI21_X1 U7873 ( .B1(alu_a_q[21]), .B2(n3839), .A(n7590), .ZN(n7578) );
  AOI222_X1 U7874 ( .A1(n7577), .A2(n7592), .B1(n3353), .B2(n7593), .C1(n7578), 
        .C2(n3352), .ZN(n7585) );
  OAI22_X1 U7875 ( .A1(n7593), .A2(n3842), .B1(n3764), .B2(n7578), .ZN(n7579)
         );
  NOR4_X1 U7876 ( .A1(n7835), .A2(n7591), .A3(n7580), .A4(n7579), .ZN(n7584)
         );
  AOI22_X1 U7877 ( .A1(alu_a_q[22]), .A2(n7802), .B1(n7801), .B2(n7807), .ZN(
        n7583) );
  AOI22_X1 U7878 ( .A1(n7796), .A2(n7679), .B1(n7808), .B2(n7581), .ZN(n7582)
         );
  OAI211_X1 U7879 ( .C1(n7585), .C2(n7584), .A(n7583), .B(n7582), .ZN(n7586)
         );
  AOI22_X1 U7880 ( .A1(n4847), .A2(n4839), .B1(n4068), .B2(n4846), .ZN(n2106)
         );
  AOI22_X1 U7881 ( .A1(n4849), .A2(n4839), .B1(n4588), .B2(n4848), .ZN(n2105)
         );
  AOI22_X1 U7882 ( .A1(n4851), .A2(n4839), .B1(n4312), .B2(n4850), .ZN(n2104)
         );
  AOI22_X1 U7883 ( .A1(n4853), .A2(n4839), .B1(n4313), .B2(n4852), .ZN(n2103)
         );
  AOI22_X1 U7884 ( .A1(n4855), .A2(n4839), .B1(n4589), .B2(n4854), .ZN(n2102)
         );
  AOI22_X1 U7885 ( .A1(n4857), .A2(n4839), .B1(n4069), .B2(n4856), .ZN(n2101)
         );
  AOI22_X1 U7886 ( .A1(n4859), .A2(n4839), .B1(n4070), .B2(n4858), .ZN(n2100)
         );
  AOI22_X1 U7887 ( .A1(n4861), .A2(n4839), .B1(n4590), .B2(n4860), .ZN(n2099)
         );
  AOI22_X1 U7888 ( .A1(n4863), .A2(n4839), .B1(n4071), .B2(n4862), .ZN(n2098)
         );
  AOI22_X1 U7889 ( .A1(n4865), .A2(n4839), .B1(n4591), .B2(n4864), .ZN(n2097)
         );
  AOI22_X1 U7890 ( .A1(n4867), .A2(n4839), .B1(n4314), .B2(n4866), .ZN(n2096)
         );
  AOI22_X1 U7891 ( .A1(n4869), .A2(n4839), .B1(n4315), .B2(n4868), .ZN(n2095)
         );
  AOI22_X1 U7892 ( .A1(n4871), .A2(n4839), .B1(n4592), .B2(n4870), .ZN(n2094)
         );
  AOI22_X1 U7893 ( .A1(n4873), .A2(n4839), .B1(n4072), .B2(n4872), .ZN(n2093)
         );
  AOI22_X1 U7894 ( .A1(n4875), .A2(n4839), .B1(n4073), .B2(n4874), .ZN(n2092)
         );
  AOI22_X1 U7895 ( .A1(n4877), .A2(n4839), .B1(n4593), .B2(n4876), .ZN(n2091)
         );
  AOI22_X1 U7896 ( .A1(n4879), .A2(n4839), .B1(n4074), .B2(n4878), .ZN(n2090)
         );
  AOI22_X1 U7897 ( .A1(n4881), .A2(n4839), .B1(n4594), .B2(n4880), .ZN(n2089)
         );
  AOI22_X1 U7898 ( .A1(n4883), .A2(n4839), .B1(n4316), .B2(n4882), .ZN(n2088)
         );
  AOI22_X1 U7899 ( .A1(n4885), .A2(n4839), .B1(n4317), .B2(n4884), .ZN(n2087)
         );
  AOI22_X1 U7900 ( .A1(n4887), .A2(n4839), .B1(n4595), .B2(n4886), .ZN(n2086)
         );
  AOI22_X1 U7901 ( .A1(n4889), .A2(n7589), .B1(n4075), .B2(n4888), .ZN(n2085)
         );
  AOI22_X1 U7902 ( .A1(n4891), .A2(n7589), .B1(n4076), .B2(n4890), .ZN(n2084)
         );
  AOI22_X1 U7903 ( .A1(n4893), .A2(n7589), .B1(n4596), .B2(n4892), .ZN(n2083)
         );
  AOI22_X1 U7904 ( .A1(n4895), .A2(n7589), .B1(n4077), .B2(n4894), .ZN(n2082)
         );
  AOI22_X1 U7905 ( .A1(n4897), .A2(n7589), .B1(n4597), .B2(n4896), .ZN(n2081)
         );
  AOI22_X1 U7906 ( .A1(n4899), .A2(n7589), .B1(n4318), .B2(n4898), .ZN(n2080)
         );
  AOI22_X1 U7907 ( .A1(n4901), .A2(n4839), .B1(n4319), .B2(n4900), .ZN(n2079)
         );
  AOI22_X1 U7908 ( .A1(n4903), .A2(n4839), .B1(n4598), .B2(n4902), .ZN(n2078)
         );
  AOI22_X1 U7909 ( .A1(n4905), .A2(n4839), .B1(n4078), .B2(n4904), .ZN(n2077)
         );
  AOI22_X1 U7910 ( .A1(n4907), .A2(n4839), .B1(n4079), .B2(n4906), .ZN(n2076)
         );
  AOI22_X1 U7911 ( .A1(n4909), .A2(n4839), .B1(n4599), .B2(n4908), .ZN(n2075)
         );
  AOI22_X1 U7912 ( .A1(alu_b_q[21]), .A2(n3766), .B1(alu_b_q[22]), .B2(n3795), 
        .ZN(n7918) );
  INV_X1 U7913 ( .A(n7630), .ZN(n7607) );
  OAI22_X1 U7914 ( .A1(n3764), .A2(n7628), .B1(n3842), .B2(n7607), .ZN(n7594)
         );
  INV_X1 U7915 ( .A(n7594), .ZN(n7595) );
  NAND2_X1 U7916 ( .A1(n3792), .A2(alu_b_q[23]), .ZN(n7643) );
  NAND2_X1 U7917 ( .A1(alu_a_q[23]), .A2(n3841), .ZN(n7923) );
  AOI22_X1 U7918 ( .A1(n7595), .A2(n7865), .B1(n7643), .B2(n7923), .ZN(n7613)
         );
  AOI22_X1 U7919 ( .A1(n7808), .A2(n7700), .B1(n7701), .B2(n7596), .ZN(n7603)
         );
  NOR4_X1 U7920 ( .A1(n7600), .A2(n7599), .A3(n7598), .A4(n7597), .ZN(n7845)
         );
  OAI22_X1 U7921 ( .A1(n7845), .A2(n7707), .B1(n7842), .B2(n7708), .ZN(n7601)
         );
  AOI21_X1 U7922 ( .B1(n7796), .B2(n7702), .A(n7601), .ZN(n7602) );
  OAI211_X1 U7923 ( .C1(n3792), .C2(n7867), .A(n7603), .B(n7602), .ZN(n7612)
         );
  AOI22_X1 U7924 ( .A1(alu_b_q[23]), .A2(n7872), .B1(n7739), .B2(n7604), .ZN(
        n7605) );
  OAI211_X1 U7925 ( .C1(n7606), .C2(n7831), .A(n7605), .B(n7797), .ZN(n7611)
         );
  AOI22_X1 U7926 ( .A1(n3352), .A2(n7628), .B1(n3353), .B2(n7607), .ZN(n7609)
         );
  NAND2_X1 U7927 ( .A1(alu_a_q[23]), .A2(alu_b_q[23]), .ZN(n7629) );
  NAND2_X1 U7928 ( .A1(n3792), .A2(n3841), .ZN(n7608) );
  AOI222_X1 U7929 ( .A1(n7609), .A2(n7629), .B1(n7609), .B2(n7788), .C1(n7629), 
        .C2(n7608), .ZN(n7610) );
  AOI22_X1 U7930 ( .A1(n4847), .A2(n3365), .B1(n4080), .B2(n4846), .ZN(n2074)
         );
  AOI22_X1 U7931 ( .A1(n4849), .A2(n3365), .B1(n4600), .B2(n4848), .ZN(n2073)
         );
  AOI22_X1 U7932 ( .A1(n4851), .A2(n3365), .B1(n4320), .B2(n4850), .ZN(n2072)
         );
  AOI22_X1 U7933 ( .A1(n4853), .A2(n3365), .B1(n4321), .B2(n4852), .ZN(n2071)
         );
  AOI22_X1 U7934 ( .A1(n4855), .A2(n3365), .B1(n4601), .B2(n4854), .ZN(n2070)
         );
  AOI22_X1 U7935 ( .A1(n4857), .A2(n3365), .B1(n4081), .B2(n4856), .ZN(n2069)
         );
  AOI22_X1 U7936 ( .A1(n4859), .A2(n3365), .B1(n4082), .B2(n4858), .ZN(n2068)
         );
  AOI22_X1 U7937 ( .A1(n4861), .A2(n3365), .B1(n4602), .B2(n4860), .ZN(n2067)
         );
  AOI22_X1 U7938 ( .A1(n4863), .A2(n3365), .B1(n4083), .B2(n4862), .ZN(n2066)
         );
  AOI22_X1 U7939 ( .A1(n4865), .A2(n3365), .B1(n4603), .B2(n4864), .ZN(n2065)
         );
  AOI22_X1 U7940 ( .A1(n4867), .A2(n3365), .B1(n4322), .B2(n4866), .ZN(n2064)
         );
  AOI22_X1 U7941 ( .A1(n4869), .A2(n3365), .B1(n4323), .B2(n4868), .ZN(n2063)
         );
  AOI22_X1 U7942 ( .A1(n4871), .A2(n7614), .B1(n4604), .B2(n4870), .ZN(n2062)
         );
  AOI22_X1 U7943 ( .A1(n4873), .A2(n7614), .B1(n4084), .B2(n4872), .ZN(n2061)
         );
  AOI22_X1 U7944 ( .A1(n4875), .A2(n3365), .B1(n4085), .B2(n4874), .ZN(n2060)
         );
  AOI22_X1 U7945 ( .A1(n4877), .A2(n3365), .B1(n4605), .B2(n4876), .ZN(n2059)
         );
  AOI22_X1 U7946 ( .A1(n4879), .A2(n3365), .B1(n4086), .B2(n4878), .ZN(n2058)
         );
  AOI22_X1 U7947 ( .A1(n4881), .A2(n3365), .B1(n4606), .B2(n4880), .ZN(n2057)
         );
  AOI22_X1 U7948 ( .A1(n4883), .A2(n3365), .B1(n4324), .B2(n4882), .ZN(n2056)
         );
  AOI22_X1 U7949 ( .A1(n4885), .A2(n3365), .B1(n4325), .B2(n4884), .ZN(n2055)
         );
  AOI22_X1 U7950 ( .A1(n4887), .A2(n3365), .B1(n4607), .B2(n4886), .ZN(n2054)
         );
  AOI22_X1 U7951 ( .A1(n4889), .A2(n3365), .B1(n4087), .B2(n4888), .ZN(n2053)
         );
  AOI22_X1 U7952 ( .A1(n4891), .A2(n3365), .B1(n4088), .B2(n4890), .ZN(n2052)
         );
  AOI22_X1 U7953 ( .A1(n4893), .A2(n3365), .B1(n4608), .B2(n4892), .ZN(n2051)
         );
  AOI22_X1 U7954 ( .A1(n4895), .A2(n3365), .B1(n4089), .B2(n4894), .ZN(n2050)
         );
  AOI22_X1 U7955 ( .A1(n4897), .A2(n3365), .B1(n4609), .B2(n4896), .ZN(n2049)
         );
  AOI22_X1 U7956 ( .A1(n4899), .A2(n3365), .B1(n4326), .B2(n4898), .ZN(n2048)
         );
  AOI22_X1 U7957 ( .A1(n4901), .A2(n3365), .B1(n4327), .B2(n4900), .ZN(n2047)
         );
  AOI22_X1 U7958 ( .A1(n4903), .A2(n3365), .B1(n4610), .B2(n4902), .ZN(n2046)
         );
  AOI22_X1 U7959 ( .A1(n4905), .A2(n3365), .B1(n4090), .B2(n4904), .ZN(n2045)
         );
  AOI22_X1 U7960 ( .A1(n4907), .A2(n3365), .B1(n4091), .B2(n4906), .ZN(n2044)
         );
  AOI22_X1 U7961 ( .A1(n4909), .A2(n3365), .B1(n4611), .B2(n4908), .ZN(n2043)
         );
  OAI22_X1 U7962 ( .A1(n7750), .A2(n7708), .B1(n3789), .B2(n7867), .ZN(n7641)
         );
  AND4_X1 U7963 ( .A1(n7618), .A2(n7617), .A3(n7616), .A4(n7615), .ZN(n7741)
         );
  NOR2_X1 U7964 ( .A1(alu_b_q[24]), .A2(n3789), .ZN(n7927) );
  INV_X1 U7965 ( .A(n7619), .ZN(n7742) );
  OAI22_X1 U7966 ( .A1(n7742), .A2(n7709), .B1(n7621), .B2(n7620), .ZN(n7622)
         );
  AOI211_X1 U7967 ( .C1(n7927), .C2(n7835), .A(n7833), .B(n7622), .ZN(n7627)
         );
  NAND2_X1 U7968 ( .A1(n3830), .A2(alu_a_q[24]), .ZN(n7623) );
  INV_X1 U7969 ( .A(n7623), .ZN(n7625) );
  OAI221_X1 U7970 ( .B1(n7625), .B2(n7624), .C1(n7623), .C2(n7856), .A(
        alu_b_q[24]), .ZN(n7626) );
  OAI211_X1 U7971 ( .C1(n7741), .C2(n7707), .A(n7627), .B(n7626), .ZN(n7640)
         );
  NAND2_X1 U7972 ( .A1(n7643), .A2(n7645), .ZN(n7631) );
  AOI22_X1 U7973 ( .A1(n3352), .A2(n7631), .B1(n3353), .B2(n7655), .ZN(n7638)
         );
  AOI22_X1 U7974 ( .A1(alu_a_q[24]), .A2(alu_b_q[24]), .B1(n3840), .B2(n3789), 
        .ZN(n7637) );
  OAI22_X1 U7975 ( .A1(n7655), .A2(n3842), .B1(n3764), .B2(n7631), .ZN(n7635)
         );
  OAI22_X1 U7976 ( .A1(n7633), .A2(n7851), .B1(n7632), .B2(n7831), .ZN(n7634)
         );
  AOI21_X1 U7977 ( .B1(n7637), .B2(n7635), .A(n7634), .ZN(n7636) );
  OAI21_X1 U7978 ( .B1(n7638), .B2(n7637), .A(n7636), .ZN(n7639) );
  AOI22_X1 U7979 ( .A1(n4847), .A2(n4840), .B1(n4092), .B2(n4846), .ZN(n2042)
         );
  AOI22_X1 U7980 ( .A1(n4849), .A2(n4840), .B1(n4612), .B2(n4848), .ZN(n2041)
         );
  AOI22_X1 U7981 ( .A1(n4851), .A2(n4840), .B1(n4328), .B2(n4850), .ZN(n2040)
         );
  AOI22_X1 U7982 ( .A1(n4853), .A2(n4840), .B1(n4329), .B2(n4852), .ZN(n2039)
         );
  AOI22_X1 U7983 ( .A1(n4855), .A2(n4840), .B1(n4613), .B2(n4854), .ZN(n2038)
         );
  AOI22_X1 U7984 ( .A1(n4857), .A2(n4840), .B1(n4093), .B2(n4856), .ZN(n2037)
         );
  AOI22_X1 U7985 ( .A1(n4859), .A2(n4840), .B1(n4094), .B2(n4858), .ZN(n2036)
         );
  AOI22_X1 U7986 ( .A1(n4861), .A2(n4840), .B1(n4614), .B2(n4860), .ZN(n2035)
         );
  AOI22_X1 U7987 ( .A1(n4863), .A2(n4840), .B1(n4095), .B2(n4862), .ZN(n2034)
         );
  AOI22_X1 U7988 ( .A1(n4865), .A2(n4840), .B1(n4615), .B2(n4864), .ZN(n2033)
         );
  AOI22_X1 U7989 ( .A1(n4867), .A2(n4840), .B1(n4330), .B2(n4866), .ZN(n2032)
         );
  AOI22_X1 U7990 ( .A1(n4869), .A2(n4840), .B1(n4331), .B2(n4868), .ZN(n2031)
         );
  AOI22_X1 U7991 ( .A1(n4871), .A2(n4840), .B1(n4616), .B2(n4870), .ZN(n2030)
         );
  AOI22_X1 U7992 ( .A1(n4873), .A2(n4840), .B1(n4096), .B2(n4872), .ZN(n2029)
         );
  AOI22_X1 U7993 ( .A1(n4875), .A2(n4840), .B1(n4097), .B2(n4874), .ZN(n2028)
         );
  AOI22_X1 U7994 ( .A1(n4877), .A2(n4840), .B1(n4617), .B2(n4876), .ZN(n2027)
         );
  AOI22_X1 U7995 ( .A1(n4879), .A2(n4840), .B1(n4098), .B2(n4878), .ZN(n2026)
         );
  AOI22_X1 U7996 ( .A1(n4881), .A2(n4840), .B1(n4618), .B2(n4880), .ZN(n2025)
         );
  AOI22_X1 U7997 ( .A1(n4883), .A2(n4840), .B1(n4332), .B2(n4882), .ZN(n2024)
         );
  AOI22_X1 U7998 ( .A1(n4885), .A2(n4840), .B1(n4333), .B2(n4884), .ZN(n2023)
         );
  AOI22_X1 U7999 ( .A1(n4887), .A2(n7642), .B1(n4619), .B2(n4886), .ZN(n2022)
         );
  AOI22_X1 U8000 ( .A1(n4889), .A2(n7642), .B1(n4099), .B2(n4888), .ZN(n2021)
         );
  AOI22_X1 U8001 ( .A1(n4891), .A2(n7642), .B1(n4100), .B2(n4890), .ZN(n2020)
         );
  AOI22_X1 U8002 ( .A1(n4893), .A2(n7642), .B1(n4620), .B2(n4892), .ZN(n2019)
         );
  AOI22_X1 U8003 ( .A1(n4895), .A2(n7642), .B1(n4101), .B2(n4894), .ZN(n2018)
         );
  AOI22_X1 U8004 ( .A1(n4897), .A2(n7642), .B1(n4621), .B2(n4896), .ZN(n2017)
         );
  AOI22_X1 U8005 ( .A1(n4899), .A2(n7642), .B1(n4334), .B2(n4898), .ZN(n2016)
         );
  AOI22_X1 U8006 ( .A1(n4901), .A2(n4840), .B1(n4335), .B2(n4900), .ZN(n2015)
         );
  AOI22_X1 U8007 ( .A1(n4903), .A2(n4840), .B1(n4622), .B2(n4902), .ZN(n2014)
         );
  AOI22_X1 U8008 ( .A1(n4905), .A2(n4840), .B1(n4102), .B2(n4904), .ZN(n2013)
         );
  AOI22_X1 U8009 ( .A1(n4907), .A2(n4840), .B1(n4103), .B2(n4906), .ZN(n2012)
         );
  AOI22_X1 U8010 ( .A1(n4909), .A2(n4840), .B1(n4623), .B2(n4908), .ZN(n2011)
         );
  OAI21_X1 U8011 ( .B1(n3840), .B2(alu_a_q[24]), .A(n7643), .ZN(n7644) );
  INV_X1 U8012 ( .A(n7644), .ZN(n7926) );
  INV_X1 U8013 ( .A(n7685), .ZN(n7661) );
  AOI221_X1 U8014 ( .B1(alu_a_q[25]), .B2(n7685), .C1(n3829), .C2(n7661), .A(
        alu_b_q[25]), .ZN(n7670) );
  OAI22_X1 U8015 ( .A1(n7647), .A2(n7831), .B1(n7646), .B2(n7851), .ZN(n7669)
         );
  NOR2_X1 U8016 ( .A1(n3829), .A2(alu_b_q[25]), .ZN(n7716) );
  AOI22_X1 U8017 ( .A1(n7835), .A2(n7716), .B1(n7796), .B2(n7648), .ZN(n7667)
         );
  NOR4_X1 U8018 ( .A1(n7652), .A2(n7651), .A3(n7650), .A4(n7649), .ZN(n7782)
         );
  INV_X1 U8019 ( .A(n7782), .ZN(n7653) );
  AOI22_X1 U8020 ( .A1(n7808), .A2(n7654), .B1(n7866), .B2(n7653), .ZN(n7666)
         );
  INV_X1 U8021 ( .A(n7655), .ZN(n7657) );
  NAND2_X1 U8022 ( .A1(alu_a_q[24]), .A2(alu_b_q[24]), .ZN(n7656) );
  AOI22_X1 U8023 ( .A1(n3789), .A2(n3840), .B1(n7657), .B2(n7656), .ZN(n7686)
         );
  OAI22_X1 U8024 ( .A1(n7781), .A2(n7708), .B1(n3829), .B2(n7867), .ZN(n7658)
         );
  AOI211_X1 U8025 ( .C1(n3353), .C2(n7659), .A(n7833), .B(n7658), .ZN(n7665)
         );
  OAI21_X1 U8026 ( .B1(n7685), .B2(n3764), .A(n7676), .ZN(n7663) );
  OAI21_X1 U8027 ( .B1(n7661), .B2(n7660), .A(n7735), .ZN(n7662) );
  OAI221_X1 U8028 ( .B1(alu_a_q[25]), .B2(n7663), .C1(n3829), .C2(n7662), .A(
        alu_b_q[25]), .ZN(n7664) );
  NAND4_X1 U8029 ( .A1(n7667), .A2(n7666), .A3(n7665), .A4(n7664), .ZN(n7668)
         );
  AOI22_X1 U8030 ( .A1(n4847), .A2(n4841), .B1(n4104), .B2(n4846), .ZN(n2010)
         );
  AOI22_X1 U8031 ( .A1(n4849), .A2(n4841), .B1(n4624), .B2(n4848), .ZN(n2009)
         );
  AOI22_X1 U8032 ( .A1(n4851), .A2(n4841), .B1(n4336), .B2(n4850), .ZN(n2008)
         );
  AOI22_X1 U8033 ( .A1(n4853), .A2(n4841), .B1(n4337), .B2(n4852), .ZN(n2007)
         );
  AOI22_X1 U8034 ( .A1(n4855), .A2(n4841), .B1(n4625), .B2(n4854), .ZN(n2006)
         );
  AOI22_X1 U8035 ( .A1(n4857), .A2(n4841), .B1(n4105), .B2(n4856), .ZN(n2005)
         );
  AOI22_X1 U8036 ( .A1(n4859), .A2(n4841), .B1(n4106), .B2(n4858), .ZN(n2004)
         );
  AOI22_X1 U8037 ( .A1(n4861), .A2(n4841), .B1(n4626), .B2(n4860), .ZN(n2003)
         );
  AOI22_X1 U8038 ( .A1(n4863), .A2(n4841), .B1(n4107), .B2(n4862), .ZN(n2002)
         );
  AOI22_X1 U8039 ( .A1(n4865), .A2(n4841), .B1(n4627), .B2(n4864), .ZN(n2001)
         );
  AOI22_X1 U8040 ( .A1(n4867), .A2(n4841), .B1(n4338), .B2(n4866), .ZN(n2000)
         );
  AOI22_X1 U8041 ( .A1(n4869), .A2(n4841), .B1(n4339), .B2(n4868), .ZN(n1999)
         );
  AOI22_X1 U8042 ( .A1(n4871), .A2(n4841), .B1(n4628), .B2(n4870), .ZN(n1998)
         );
  AOI22_X1 U8043 ( .A1(n4873), .A2(n4841), .B1(n4108), .B2(n4872), .ZN(n1997)
         );
  AOI22_X1 U8044 ( .A1(n4875), .A2(n4841), .B1(n4109), .B2(n4874), .ZN(n1996)
         );
  AOI22_X1 U8045 ( .A1(n4877), .A2(n4841), .B1(n4629), .B2(n4876), .ZN(n1995)
         );
  AOI22_X1 U8046 ( .A1(n4879), .A2(n4841), .B1(n4110), .B2(n4878), .ZN(n1994)
         );
  AOI22_X1 U8047 ( .A1(n4881), .A2(n4841), .B1(n4630), .B2(n4880), .ZN(n1993)
         );
  AOI22_X1 U8048 ( .A1(n4883), .A2(n4841), .B1(n4340), .B2(n4882), .ZN(n1992)
         );
  AOI22_X1 U8049 ( .A1(n4885), .A2(n4841), .B1(n4341), .B2(n4884), .ZN(n1991)
         );
  AOI22_X1 U8050 ( .A1(n4887), .A2(n4841), .B1(n4631), .B2(n4886), .ZN(n1990)
         );
  AOI22_X1 U8051 ( .A1(n4889), .A2(n7671), .B1(n4111), .B2(n4888), .ZN(n1989)
         );
  AOI22_X1 U8052 ( .A1(n4891), .A2(n7671), .B1(n4112), .B2(n4890), .ZN(n1988)
         );
  AOI22_X1 U8053 ( .A1(n4893), .A2(n7671), .B1(n4632), .B2(n4892), .ZN(n1987)
         );
  AOI22_X1 U8054 ( .A1(n4895), .A2(n7671), .B1(n4113), .B2(n4894), .ZN(n1986)
         );
  AOI22_X1 U8055 ( .A1(n4897), .A2(n7671), .B1(n4633), .B2(n4896), .ZN(n1985)
         );
  AOI22_X1 U8056 ( .A1(n4899), .A2(n7671), .B1(n4342), .B2(n4898), .ZN(n1984)
         );
  AOI22_X1 U8057 ( .A1(n4901), .A2(n4841), .B1(n4343), .B2(n4900), .ZN(n1983)
         );
  AOI22_X1 U8058 ( .A1(n4903), .A2(n4841), .B1(n4634), .B2(n4902), .ZN(n1982)
         );
  AOI22_X1 U8059 ( .A1(n4905), .A2(n4841), .B1(n4114), .B2(n4904), .ZN(n1981)
         );
  AOI22_X1 U8060 ( .A1(n4907), .A2(n4841), .B1(n4115), .B2(n4906), .ZN(n1980)
         );
  AOI22_X1 U8061 ( .A1(n4909), .A2(n4841), .B1(n4635), .B2(n4908), .ZN(n1979)
         );
  NOR3_X1 U8062 ( .A1(n157), .A2(n3832), .A3(n3783), .ZN(n7677) );
  AOI22_X1 U8063 ( .A1(n7856), .A2(n7677), .B1(n7801), .B2(n7795), .ZN(n7682)
         );
  NAND4_X1 U8064 ( .A1(n7675), .A2(n7674), .A3(n7673), .A4(n7672), .ZN(n7800)
         );
  AOI22_X1 U8065 ( .A1(n7796), .A2(n7807), .B1(n7866), .B2(n7800), .ZN(n7681)
         );
  AOI211_X1 U8066 ( .C1(n157), .C2(n3783), .A(n7677), .B(n7676), .ZN(n7678) );
  NAND2_X1 U8067 ( .A1(n3832), .A2(n3783), .ZN(n7714) );
  AOI22_X1 U8068 ( .A1(n7808), .A2(n7679), .B1(n7678), .B2(n7714), .ZN(n7680)
         );
  NAND4_X1 U8069 ( .A1(n7682), .A2(n7681), .A3(n7680), .A4(n7797), .ZN(n7695)
         );
  OAI22_X1 U8070 ( .A1(n7684), .A2(n7851), .B1(n7683), .B2(n7831), .ZN(n7694)
         );
  NOR2_X1 U8071 ( .A1(n7716), .A2(n7718), .ZN(n7687) );
  FA_X1 U8072 ( .A(alu_b_q[25]), .B(alu_a_q[25]), .CI(n7686), .CO(n7715), .S(
        n7659) );
  AOI22_X1 U8073 ( .A1(n3352), .A2(n7687), .B1(n7715), .B2(n3353), .ZN(n7692)
         );
  OAI21_X1 U8074 ( .B1(n7692), .B2(n3783), .A(n7867), .ZN(n7690) );
  OAI22_X1 U8075 ( .A1(n7715), .A2(n3842), .B1(n7687), .B2(n3764), .ZN(n7689)
         );
  XOR2_X1 U8076 ( .A(n3832), .B(n3783), .Z(n7688) );
  AOI22_X1 U8077 ( .A1(alu_a_q[26]), .A2(n7690), .B1(n7689), .B2(n7688), .ZN(
        n7691) );
  OAI21_X1 U8078 ( .B1(n7692), .B2(n7714), .A(n7691), .ZN(n7693) );
  AOI22_X1 U8079 ( .A1(n7954), .A2(n4842), .B1(n4116), .B2(n4846), .ZN(n1978)
         );
  AOI22_X1 U8080 ( .A1(n7955), .A2(n4842), .B1(n4636), .B2(n4848), .ZN(n1977)
         );
  AOI22_X1 U8081 ( .A1(n7956), .A2(n4842), .B1(n4344), .B2(n4850), .ZN(n1976)
         );
  AOI22_X1 U8082 ( .A1(n7957), .A2(n4842), .B1(n4345), .B2(n4852), .ZN(n1975)
         );
  AOI22_X1 U8083 ( .A1(n7958), .A2(n4842), .B1(n4637), .B2(n4854), .ZN(n1974)
         );
  AOI22_X1 U8084 ( .A1(n7959), .A2(n4842), .B1(n4117), .B2(n4856), .ZN(n1973)
         );
  AOI22_X1 U8085 ( .A1(n7960), .A2(n4842), .B1(n4118), .B2(n4858), .ZN(n1972)
         );
  AOI22_X1 U8086 ( .A1(n7961), .A2(n4842), .B1(n4638), .B2(n4860), .ZN(n1971)
         );
  AOI22_X1 U8087 ( .A1(n7962), .A2(n4842), .B1(n4119), .B2(n4862), .ZN(n1970)
         );
  AOI22_X1 U8088 ( .A1(n7963), .A2(n4842), .B1(n4639), .B2(n4864), .ZN(n1969)
         );
  AOI22_X1 U8089 ( .A1(n7964), .A2(n4842), .B1(n4346), .B2(n4866), .ZN(n1968)
         );
  AOI22_X1 U8090 ( .A1(n7965), .A2(n4842), .B1(n4347), .B2(n4868), .ZN(n1967)
         );
  AOI22_X1 U8091 ( .A1(n7966), .A2(n4842), .B1(n4640), .B2(n4870), .ZN(n1966)
         );
  AOI22_X1 U8092 ( .A1(n7967), .A2(n4842), .B1(n4120), .B2(n4872), .ZN(n1965)
         );
  AOI22_X1 U8093 ( .A1(n7968), .A2(n4842), .B1(n4121), .B2(n4874), .ZN(n1964)
         );
  AOI22_X1 U8094 ( .A1(n7969), .A2(n4842), .B1(n4641), .B2(n4876), .ZN(n1963)
         );
  AOI22_X1 U8095 ( .A1(n7970), .A2(n4842), .B1(n4122), .B2(n4878), .ZN(n1962)
         );
  AOI22_X1 U8096 ( .A1(n7971), .A2(n4842), .B1(n4642), .B2(n4880), .ZN(n1961)
         );
  AOI22_X1 U8097 ( .A1(n7972), .A2(n4842), .B1(n4348), .B2(n4882), .ZN(n1960)
         );
  AOI22_X1 U8098 ( .A1(n7973), .A2(n4842), .B1(n4349), .B2(n4884), .ZN(n1959)
         );
  AOI22_X1 U8099 ( .A1(n4887), .A2(n7696), .B1(n4643), .B2(n4886), .ZN(n1958)
         );
  AOI22_X1 U8100 ( .A1(n4889), .A2(n7696), .B1(n4123), .B2(n4888), .ZN(n1957)
         );
  AOI22_X1 U8101 ( .A1(n4891), .A2(n7696), .B1(n4124), .B2(n4890), .ZN(n1956)
         );
  AOI22_X1 U8102 ( .A1(n4893), .A2(n7696), .B1(n4644), .B2(n4892), .ZN(n1955)
         );
  AOI22_X1 U8103 ( .A1(n4895), .A2(n7696), .B1(n4125), .B2(n4894), .ZN(n1954)
         );
  AOI22_X1 U8104 ( .A1(n4897), .A2(n7696), .B1(n4645), .B2(n4896), .ZN(n1953)
         );
  AOI22_X1 U8105 ( .A1(n4899), .A2(n7696), .B1(n4350), .B2(n4898), .ZN(n1952)
         );
  AOI22_X1 U8106 ( .A1(n7981), .A2(n4842), .B1(n4351), .B2(n4900), .ZN(n1951)
         );
  AOI22_X1 U8107 ( .A1(n7982), .A2(n4842), .B1(n4646), .B2(n4902), .ZN(n1950)
         );
  AOI22_X1 U8108 ( .A1(n7983), .A2(n4842), .B1(n4126), .B2(n4904), .ZN(n1949)
         );
  AOI22_X1 U8109 ( .A1(n7984), .A2(n4842), .B1(n4127), .B2(n4906), .ZN(n1948)
         );
  AOI22_X1 U8110 ( .A1(n7985), .A2(n4842), .B1(n4647), .B2(n4908), .ZN(n1947)
         );
  AOI22_X1 U8111 ( .A1(n7699), .A2(n7698), .B1(n7739), .B2(n7697), .ZN(n7727)
         );
  AOI22_X1 U8112 ( .A1(n7808), .A2(n7702), .B1(n7701), .B2(n7700), .ZN(n7726)
         );
  NAND2_X1 U8113 ( .A1(alu_a_q[27]), .A2(alu_b_q[27]), .ZN(n7732) );
  OAI22_X1 U8114 ( .A1(n3784), .A2(n7867), .B1(n7732), .B2(n7788), .ZN(n7712)
         );
  NOR4_X1 U8115 ( .A1(n7706), .A2(n7705), .A3(n7704), .A4(n7703), .ZN(n7844)
         );
  OAI22_X1 U8116 ( .A1(n7845), .A2(n7708), .B1(n7844), .B2(n7707), .ZN(n7711)
         );
  OAI22_X1 U8117 ( .A1(n7842), .A2(n7709), .B1(n3843), .B2(n7734), .ZN(n7710)
         );
  NOR4_X1 U8118 ( .A1(n7833), .A2(n7712), .A3(n7711), .A4(n7710), .ZN(n7725)
         );
  NOR2_X1 U8119 ( .A1(n3784), .A2(alu_b_q[27]), .ZN(n7765) );
  AOI21_X1 U8120 ( .B1(n3784), .B2(alu_b_q[27]), .A(n7765), .ZN(n7713) );
  INV_X1 U8121 ( .A(n7713), .ZN(n7723) );
  NOR2_X1 U8122 ( .A1(n3783), .A2(alu_a_q[26]), .ZN(n7729) );
  AOI21_X1 U8123 ( .B1(n3783), .B2(alu_a_q[26]), .A(n7716), .ZN(n7717) );
  INV_X1 U8124 ( .A(n7717), .ZN(n7889) );
  NOR2_X1 U8125 ( .A1(n7729), .A2(n7731), .ZN(n7719) );
  OAI22_X1 U8126 ( .A1(n7733), .A2(n3842), .B1(n7719), .B2(n3764), .ZN(n7722)
         );
  AOI22_X1 U8127 ( .A1(n3352), .A2(n7719), .B1(n7733), .B2(n3353), .ZN(n7720)
         );
  NAND3_X1 U8128 ( .A1(n7723), .A2(n7720), .A3(n7865), .ZN(n7721) );
  OAI21_X1 U8129 ( .B1(n7723), .B2(n7722), .A(n7721), .ZN(n7724) );
  AOI22_X1 U8130 ( .A1(n7954), .A2(n7728), .B1(n4128), .B2(n4846), .ZN(n1946)
         );
  AOI22_X1 U8131 ( .A1(n7955), .A2(n7728), .B1(n4648), .B2(n4848), .ZN(n1945)
         );
  AOI22_X1 U8132 ( .A1(n7956), .A2(n7728), .B1(n4352), .B2(n4850), .ZN(n1944)
         );
  AOI22_X1 U8133 ( .A1(n7957), .A2(n7728), .B1(n4353), .B2(n4852), .ZN(n1943)
         );
  AOI22_X1 U8134 ( .A1(n7958), .A2(n7728), .B1(n4649), .B2(n4854), .ZN(n1942)
         );
  AOI22_X1 U8135 ( .A1(n7959), .A2(n7728), .B1(n4129), .B2(n4856), .ZN(n1941)
         );
  AOI22_X1 U8136 ( .A1(n7960), .A2(n7728), .B1(n4130), .B2(n4858), .ZN(n1940)
         );
  AOI22_X1 U8137 ( .A1(n7961), .A2(n7728), .B1(n4650), .B2(n4860), .ZN(n1939)
         );
  AOI22_X1 U8138 ( .A1(n7962), .A2(n7728), .B1(n4131), .B2(n4862), .ZN(n1938)
         );
  AOI22_X1 U8139 ( .A1(n7963), .A2(n7728), .B1(n4651), .B2(n4864), .ZN(n1937)
         );
  AOI22_X1 U8140 ( .A1(n7964), .A2(n7728), .B1(n4354), .B2(n4866), .ZN(n1936)
         );
  AOI22_X1 U8141 ( .A1(n7965), .A2(n7728), .B1(n4355), .B2(n4868), .ZN(n1935)
         );
  AOI22_X1 U8142 ( .A1(n4871), .A2(n7728), .B1(n4652), .B2(n4870), .ZN(n1934)
         );
  AOI22_X1 U8143 ( .A1(n4873), .A2(n7728), .B1(n4132), .B2(n4872), .ZN(n1933)
         );
  AOI22_X1 U8144 ( .A1(n4875), .A2(n7728), .B1(n4133), .B2(n4874), .ZN(n1932)
         );
  AOI22_X1 U8145 ( .A1(n4877), .A2(n7728), .B1(n4653), .B2(n4876), .ZN(n1931)
         );
  AOI22_X1 U8146 ( .A1(n4879), .A2(n7728), .B1(n4134), .B2(n4878), .ZN(n1930)
         );
  AOI22_X1 U8147 ( .A1(n4881), .A2(n7728), .B1(n4654), .B2(n4880), .ZN(n1929)
         );
  AOI22_X1 U8148 ( .A1(n4883), .A2(n7728), .B1(n4356), .B2(n4882), .ZN(n1928)
         );
  AOI22_X1 U8149 ( .A1(n4885), .A2(n7728), .B1(n4357), .B2(n4884), .ZN(n1927)
         );
  AOI22_X1 U8150 ( .A1(n4887), .A2(n7728), .B1(n4655), .B2(n4886), .ZN(n1926)
         );
  AOI22_X1 U8151 ( .A1(n4889), .A2(n7728), .B1(n4135), .B2(n4888), .ZN(n1925)
         );
  AOI22_X1 U8152 ( .A1(n4891), .A2(n7728), .B1(n4136), .B2(n4890), .ZN(n1924)
         );
  AOI22_X1 U8153 ( .A1(n4893), .A2(n7728), .B1(n4656), .B2(n4892), .ZN(n1923)
         );
  AOI22_X1 U8154 ( .A1(n4895), .A2(n7728), .B1(n4137), .B2(n4894), .ZN(n1922)
         );
  AOI22_X1 U8155 ( .A1(n4897), .A2(n7728), .B1(n4657), .B2(n4896), .ZN(n1921)
         );
  AOI22_X1 U8156 ( .A1(n4899), .A2(n7728), .B1(n4358), .B2(n4898), .ZN(n1920)
         );
  AOI22_X1 U8157 ( .A1(n7981), .A2(n7728), .B1(n4359), .B2(n4900), .ZN(n1919)
         );
  AOI22_X1 U8158 ( .A1(n7982), .A2(n7728), .B1(n4658), .B2(n4902), .ZN(n1918)
         );
  AOI22_X1 U8159 ( .A1(n4905), .A2(n7728), .B1(n4138), .B2(n4904), .ZN(n1917)
         );
  AOI22_X1 U8160 ( .A1(n7984), .A2(n7728), .B1(n4139), .B2(n4906), .ZN(n1916)
         );
  AOI22_X1 U8161 ( .A1(n4909), .A2(n7728), .B1(n4659), .B2(n4908), .ZN(n1915)
         );
  AOI21_X1 U8162 ( .B1(n3784), .B2(alu_b_q[27]), .A(n7729), .ZN(n7730) );
  INV_X1 U8163 ( .A(n7730), .ZN(n7930) );
  NOR2_X1 U8164 ( .A1(n7765), .A2(n7767), .ZN(n7757) );
  AOI22_X1 U8165 ( .A1(n3352), .A2(n7757), .B1(n7769), .B2(n3353), .ZN(n7756)
         );
  AOI22_X1 U8166 ( .A1(n7735), .A2(n7756), .B1(n3790), .B2(n7734), .ZN(n7763)
         );
  NAND2_X1 U8167 ( .A1(n3790), .A2(n3834), .ZN(n7768) );
  OAI22_X1 U8168 ( .A1(n3790), .A2(n7867), .B1(n7831), .B2(n7736), .ZN(n7737)
         );
  AOI211_X1 U8169 ( .C1(n7739), .C2(n7738), .A(n7833), .B(n7737), .ZN(n7755)
         );
  INV_X1 U8170 ( .A(n7740), .ZN(n7843) );
  OAI22_X1 U8171 ( .A1(n7742), .A2(n7877), .B1(n7741), .B2(n7843), .ZN(n7753)
         );
  NAND2_X1 U8172 ( .A1(alu_a_q[28]), .A2(n7743), .ZN(n7746) );
  AND4_X1 U8173 ( .A1(n7747), .A2(n7746), .A3(n7745), .A4(n7744), .ZN(n7751)
         );
  INV_X1 U8174 ( .A(n7748), .ZN(n7840) );
  INV_X1 U8175 ( .A(n7749), .ZN(n7879) );
  OAI22_X1 U8176 ( .A1(n7751), .A2(n7840), .B1(n7750), .B2(n7879), .ZN(n7752)
         );
  OAI21_X1 U8177 ( .B1(n7753), .B2(n7752), .A(n7846), .ZN(n7754) );
  OAI211_X1 U8178 ( .C1(n7756), .C2(n7768), .A(n7755), .B(n7754), .ZN(n7762)
         );
  NOR2_X1 U8179 ( .A1(n3834), .A2(alu_a_q[28]), .ZN(n7928) );
  INV_X1 U8180 ( .A(n7928), .ZN(n7766) );
  NAND2_X1 U8181 ( .A1(alu_a_q[28]), .A2(n3834), .ZN(n7760) );
  OAI22_X1 U8182 ( .A1(n7769), .A2(n3842), .B1(n7757), .B2(n3764), .ZN(n7758)
         );
  NOR2_X1 U8183 ( .A1(n7835), .A2(n7758), .ZN(n7759) );
  AOI21_X1 U8184 ( .B1(n7766), .B2(n7760), .A(n7759), .ZN(n7761) );
  AOI22_X1 U8185 ( .A1(n7954), .A2(n4843), .B1(n4140), .B2(n4846), .ZN(n1914)
         );
  AOI22_X1 U8186 ( .A1(n7955), .A2(n4843), .B1(n4660), .B2(n4848), .ZN(n1913)
         );
  AOI22_X1 U8187 ( .A1(n7956), .A2(n4843), .B1(n4360), .B2(n4850), .ZN(n1912)
         );
  AOI22_X1 U8188 ( .A1(n7957), .A2(n4843), .B1(n4361), .B2(n4852), .ZN(n1911)
         );
  AOI22_X1 U8189 ( .A1(n7958), .A2(n4843), .B1(n4661), .B2(n4854), .ZN(n1910)
         );
  AOI22_X1 U8190 ( .A1(n7959), .A2(n4843), .B1(n4141), .B2(n4856), .ZN(n1909)
         );
  AOI22_X1 U8191 ( .A1(n7960), .A2(n4843), .B1(n4142), .B2(n4858), .ZN(n1908)
         );
  AOI22_X1 U8192 ( .A1(n7961), .A2(n4843), .B1(n4662), .B2(n4860), .ZN(n1907)
         );
  AOI22_X1 U8193 ( .A1(n7962), .A2(n4843), .B1(n4143), .B2(n4862), .ZN(n1906)
         );
  AOI22_X1 U8194 ( .A1(n7963), .A2(n4843), .B1(n4663), .B2(n4864), .ZN(n1905)
         );
  AOI22_X1 U8195 ( .A1(n7964), .A2(n4843), .B1(n4362), .B2(n4866), .ZN(n1904)
         );
  AOI22_X1 U8196 ( .A1(n7965), .A2(n4843), .B1(n4363), .B2(n4868), .ZN(n1903)
         );
  AOI22_X1 U8197 ( .A1(n7966), .A2(n4843), .B1(n4664), .B2(n4870), .ZN(n1902)
         );
  AOI22_X1 U8198 ( .A1(n7967), .A2(n4843), .B1(n4144), .B2(n4872), .ZN(n1901)
         );
  AOI22_X1 U8199 ( .A1(n7968), .A2(n4843), .B1(n4145), .B2(n4874), .ZN(n1900)
         );
  AOI22_X1 U8200 ( .A1(n7969), .A2(n4843), .B1(n4665), .B2(n4876), .ZN(n1899)
         );
  AOI22_X1 U8201 ( .A1(n7970), .A2(n4843), .B1(n4146), .B2(n4878), .ZN(n1898)
         );
  AOI22_X1 U8202 ( .A1(n7971), .A2(n4843), .B1(n4666), .B2(n4880), .ZN(n1897)
         );
  AOI22_X1 U8203 ( .A1(n7972), .A2(n4843), .B1(n4364), .B2(n4882), .ZN(n1896)
         );
  AOI22_X1 U8204 ( .A1(n7973), .A2(n4843), .B1(n4365), .B2(n4884), .ZN(n1895)
         );
  AOI22_X1 U8205 ( .A1(n7974), .A2(n4843), .B1(n4667), .B2(n4886), .ZN(n1894)
         );
  AOI22_X1 U8206 ( .A1(n7975), .A2(n7764), .B1(n4147), .B2(n4888), .ZN(n1893)
         );
  AOI22_X1 U8207 ( .A1(n7976), .A2(n7764), .B1(n4148), .B2(n4890), .ZN(n1892)
         );
  AOI22_X1 U8208 ( .A1(n7977), .A2(n7764), .B1(n4668), .B2(n4892), .ZN(n1891)
         );
  AOI22_X1 U8209 ( .A1(n4895), .A2(n7764), .B1(n4149), .B2(n4894), .ZN(n1890)
         );
  AOI22_X1 U8210 ( .A1(n4897), .A2(n7764), .B1(n4669), .B2(n4896), .ZN(n1889)
         );
  AOI22_X1 U8211 ( .A1(n4899), .A2(n7764), .B1(n4366), .B2(n4898), .ZN(n1888)
         );
  AOI22_X1 U8212 ( .A1(n7981), .A2(n4843), .B1(n4367), .B2(n4900), .ZN(n1887)
         );
  AOI22_X1 U8213 ( .A1(n7982), .A2(n4843), .B1(n4670), .B2(n4902), .ZN(n1886)
         );
  AOI22_X1 U8214 ( .A1(n7983), .A2(n4843), .B1(n4150), .B2(n4904), .ZN(n1885)
         );
  AOI22_X1 U8215 ( .A1(n7984), .A2(n4843), .B1(n4151), .B2(n4906), .ZN(n1884)
         );
  AOI22_X1 U8216 ( .A1(n7985), .A2(n4843), .B1(n4671), .B2(n4908), .ZN(n1883)
         );
  AOI21_X1 U8217 ( .B1(n3834), .B2(alu_a_q[28]), .A(n7765), .ZN(n7931) );
  INV_X1 U8218 ( .A(n7931), .ZN(n7888) );
  AOI22_X1 U8219 ( .A1(alu_a_q[28]), .A2(alu_b_q[28]), .B1(n7769), .B2(n7768), 
        .ZN(n7818) );
  INV_X1 U8220 ( .A(n7818), .ZN(n7787) );
  OAI22_X1 U8221 ( .A1(n3764), .A2(n7813), .B1(n7787), .B2(n3842), .ZN(n7770)
         );
  NAND2_X1 U8222 ( .A1(n3836), .A2(alu_a_q[29]), .ZN(n7828) );
  INV_X1 U8223 ( .A(n7828), .ZN(n7814) );
  NOR2_X1 U8224 ( .A1(alu_a_q[29]), .A2(n3836), .ZN(n7929) );
  OAI22_X1 U8225 ( .A1(n7770), .A2(n7835), .B1(n7814), .B2(n7929), .ZN(n7771)
         );
  INV_X1 U8226 ( .A(n7771), .ZN(n7793) );
  AOI22_X1 U8227 ( .A1(alu_a_q[29]), .A2(n7802), .B1(alu_b_q[29]), .B2(n7872), 
        .ZN(n7772) );
  OAI211_X1 U8228 ( .C1(n7773), .C2(n7851), .A(n7772), .B(n7797), .ZN(n7792)
         );
  NOR2_X1 U8229 ( .A1(n3797), .A2(n7774), .ZN(n7778) );
  NOR4_X1 U8230 ( .A1(n7778), .A2(n7777), .A3(n7776), .A4(n7775), .ZN(n7780)
         );
  OAI22_X1 U8231 ( .A1(n7780), .A2(n7840), .B1(n7779), .B2(n7877), .ZN(n7784)
         );
  OAI22_X1 U8232 ( .A1(n7782), .A2(n7843), .B1(n7781), .B2(n7879), .ZN(n7783)
         );
  OAI21_X1 U8233 ( .B1(n7784), .B2(n7783), .A(n7846), .ZN(n7785) );
  OAI21_X1 U8234 ( .B1(n7831), .B2(n7786), .A(n7785), .ZN(n7791) );
  AOI22_X1 U8235 ( .A1(n3352), .A2(n7813), .B1(n3353), .B2(n7787), .ZN(n7789)
         );
  NAND2_X1 U8236 ( .A1(alu_a_q[29]), .A2(alu_b_q[29]), .ZN(n7817) );
  NAND2_X1 U8237 ( .A1(n3797), .A2(n3836), .ZN(n7815) );
  AOI222_X1 U8238 ( .A1(n7789), .A2(n7817), .B1(n7789), .B2(n7788), .C1(n7817), 
        .C2(n7815), .ZN(n7790) );
  AOI22_X1 U8239 ( .A1(n4847), .A2(n3364), .B1(n4152), .B2(n4846), .ZN(n1882)
         );
  AOI22_X1 U8240 ( .A1(n4849), .A2(n3364), .B1(n4672), .B2(n4848), .ZN(n1881)
         );
  AOI22_X1 U8241 ( .A1(n4851), .A2(n3364), .B1(n4368), .B2(n4850), .ZN(n1880)
         );
  AOI22_X1 U8242 ( .A1(n4853), .A2(n3364), .B1(n4369), .B2(n4852), .ZN(n1879)
         );
  AOI22_X1 U8243 ( .A1(n4855), .A2(n3364), .B1(n4673), .B2(n4854), .ZN(n1878)
         );
  AOI22_X1 U8244 ( .A1(n4857), .A2(n3364), .B1(n4153), .B2(n4856), .ZN(n1877)
         );
  AOI22_X1 U8245 ( .A1(n4859), .A2(n3364), .B1(n4154), .B2(n4858), .ZN(n1876)
         );
  AOI22_X1 U8246 ( .A1(n4861), .A2(n3364), .B1(n4674), .B2(n4860), .ZN(n1875)
         );
  AOI22_X1 U8247 ( .A1(n4863), .A2(n3364), .B1(n4155), .B2(n4862), .ZN(n1874)
         );
  AOI22_X1 U8248 ( .A1(n4865), .A2(n3364), .B1(n4675), .B2(n4864), .ZN(n1873)
         );
  AOI22_X1 U8249 ( .A1(n4867), .A2(n3364), .B1(n4370), .B2(n4866), .ZN(n1872)
         );
  AOI22_X1 U8250 ( .A1(n4869), .A2(n3364), .B1(n4371), .B2(n4868), .ZN(n1871)
         );
  AOI22_X1 U8251 ( .A1(n7966), .A2(n3364), .B1(n4676), .B2(n4870), .ZN(n1870)
         );
  AOI22_X1 U8252 ( .A1(n7967), .A2(n3364), .B1(n4156), .B2(n4872), .ZN(n1869)
         );
  AOI22_X1 U8253 ( .A1(n7968), .A2(n3364), .B1(n4157), .B2(n4874), .ZN(n1868)
         );
  AOI22_X1 U8254 ( .A1(n7969), .A2(n3364), .B1(n4677), .B2(n4876), .ZN(n1867)
         );
  AOI22_X1 U8255 ( .A1(n4879), .A2(n3364), .B1(n4158), .B2(n4878), .ZN(n1866)
         );
  AOI22_X1 U8256 ( .A1(n4881), .A2(n3364), .B1(n4678), .B2(n4880), .ZN(n1865)
         );
  AOI22_X1 U8257 ( .A1(n4883), .A2(n3364), .B1(n4372), .B2(n4882), .ZN(n1864)
         );
  AOI22_X1 U8258 ( .A1(n4885), .A2(n3364), .B1(n4373), .B2(n4884), .ZN(n1863)
         );
  AOI22_X1 U8259 ( .A1(n7974), .A2(n3364), .B1(n4679), .B2(n4886), .ZN(n1862)
         );
  AOI22_X1 U8260 ( .A1(n7975), .A2(n3364), .B1(n4159), .B2(n4888), .ZN(n1861)
         );
  AOI22_X1 U8261 ( .A1(n7976), .A2(n3364), .B1(n4160), .B2(n4890), .ZN(n1860)
         );
  AOI22_X1 U8262 ( .A1(n7977), .A2(n3364), .B1(n4680), .B2(n4892), .ZN(n1859)
         );
  AOI22_X1 U8263 ( .A1(n7978), .A2(n3364), .B1(n4161), .B2(n4894), .ZN(n1858)
         );
  AOI22_X1 U8264 ( .A1(n7979), .A2(n3364), .B1(n4681), .B2(n4896), .ZN(n1857)
         );
  AOI22_X1 U8265 ( .A1(n7980), .A2(n3364), .B1(n4374), .B2(n4898), .ZN(n1856)
         );
  AOI22_X1 U8266 ( .A1(n4901), .A2(n3364), .B1(n4375), .B2(n4900), .ZN(n1855)
         );
  AOI22_X1 U8267 ( .A1(n4903), .A2(n3364), .B1(n4682), .B2(n4902), .ZN(n1854)
         );
  AOI22_X1 U8268 ( .A1(n4905), .A2(n3364), .B1(n4162), .B2(n4904), .ZN(n1853)
         );
  AOI22_X1 U8269 ( .A1(n4907), .A2(n3364), .B1(n4163), .B2(n4906), .ZN(n1852)
         );
  AOI22_X1 U8270 ( .A1(n4909), .A2(n3364), .B1(n4683), .B2(n4908), .ZN(n1851)
         );
  AOI22_X1 U8271 ( .A1(alu_b_q[30]), .A2(n7872), .B1(n7796), .B2(n7795), .ZN(
        n7798) );
  OAI211_X1 U8272 ( .C1(n7831), .C2(n7799), .A(n7798), .B(n7797), .ZN(n7826)
         );
  AOI22_X1 U8273 ( .A1(alu_a_q[30]), .A2(n7802), .B1(n7801), .B2(n7800), .ZN(
        n7811) );
  NAND4_X1 U8274 ( .A1(n7806), .A2(n7805), .A3(n7804), .A4(n7803), .ZN(n7809)
         );
  AOI22_X1 U8275 ( .A1(n7866), .A2(n7809), .B1(n7808), .B2(n7807), .ZN(n7810)
         );
  OAI211_X1 U8276 ( .C1(n7812), .C2(n7851), .A(n7811), .B(n7810), .ZN(n7825)
         );
  NOR2_X1 U8277 ( .A1(n7814), .A2(n7829), .ZN(n7819) );
  INV_X1 U8278 ( .A(n7815), .ZN(n7816) );
  AOI222_X1 U8279 ( .A1(n3352), .A2(n7819), .B1(n7853), .B2(n3353), .C1(
        alu_b_q[30]), .C2(n7871), .ZN(n7823) );
  NAND2_X1 U8280 ( .A1(alu_b_q[30]), .A2(n3833), .ZN(n7933) );
  OAI21_X1 U8281 ( .B1(alu_b_q[30]), .B2(n3833), .A(n7933), .ZN(n7822) );
  OAI22_X1 U8282 ( .A1(n7819), .A2(n3764), .B1(n7853), .B2(n3842), .ZN(n7820)
         );
  OAI21_X1 U8283 ( .B1(n7820), .B2(n7835), .A(n7822), .ZN(n7821) );
  OAI21_X1 U8284 ( .B1(n7823), .B2(n7822), .A(n7821), .ZN(n7824) );
  AOI22_X1 U8285 ( .A1(n7954), .A2(n4844), .B1(n4164), .B2(n4846), .ZN(n1850)
         );
  AOI22_X1 U8286 ( .A1(n7955), .A2(n4844), .B1(n4684), .B2(n4848), .ZN(n1849)
         );
  AOI22_X1 U8287 ( .A1(n7956), .A2(n4844), .B1(n4376), .B2(n4850), .ZN(n1848)
         );
  AOI22_X1 U8288 ( .A1(n7957), .A2(n4844), .B1(n4377), .B2(n4852), .ZN(n1847)
         );
  AOI22_X1 U8289 ( .A1(n7958), .A2(n4844), .B1(n4685), .B2(n4854), .ZN(n1846)
         );
  AOI22_X1 U8290 ( .A1(n7959), .A2(n4844), .B1(n4165), .B2(n4856), .ZN(n1845)
         );
  AOI22_X1 U8291 ( .A1(n7960), .A2(n4844), .B1(n4166), .B2(n4858), .ZN(n1844)
         );
  AOI22_X1 U8292 ( .A1(n7961), .A2(n4844), .B1(n4686), .B2(n4860), .ZN(n1843)
         );
  AOI22_X1 U8293 ( .A1(n7962), .A2(n4844), .B1(n4167), .B2(n4862), .ZN(n1842)
         );
  AOI22_X1 U8294 ( .A1(n7963), .A2(n4844), .B1(n4687), .B2(n4864), .ZN(n1841)
         );
  AOI22_X1 U8295 ( .A1(n7964), .A2(n4844), .B1(n4378), .B2(n4866), .ZN(n1840)
         );
  AOI22_X1 U8296 ( .A1(n7965), .A2(n4844), .B1(n4379), .B2(n4868), .ZN(n1839)
         );
  AOI22_X1 U8297 ( .A1(n7966), .A2(n4844), .B1(n4688), .B2(n4870), .ZN(n1838)
         );
  AOI22_X1 U8298 ( .A1(n7967), .A2(n4844), .B1(n4168), .B2(n4872), .ZN(n1837)
         );
  AOI22_X1 U8299 ( .A1(n7968), .A2(n4844), .B1(n4169), .B2(n4874), .ZN(n1836)
         );
  AOI22_X1 U8300 ( .A1(n7969), .A2(n4844), .B1(n4689), .B2(n4876), .ZN(n1835)
         );
  AOI22_X1 U8301 ( .A1(n7970), .A2(n4844), .B1(n4170), .B2(n4878), .ZN(n1834)
         );
  AOI22_X1 U8302 ( .A1(n7971), .A2(n4844), .B1(n4690), .B2(n4880), .ZN(n1833)
         );
  AOI22_X1 U8303 ( .A1(n7972), .A2(n4844), .B1(n4380), .B2(n4882), .ZN(n1832)
         );
  AOI22_X1 U8304 ( .A1(n7973), .A2(n4844), .B1(n4381), .B2(n4884), .ZN(n1831)
         );
  AOI22_X1 U8305 ( .A1(n7974), .A2(n7827), .B1(n4691), .B2(n4886), .ZN(n1830)
         );
  AOI22_X1 U8306 ( .A1(n7975), .A2(n7827), .B1(n4171), .B2(n4888), .ZN(n1829)
         );
  AOI22_X1 U8307 ( .A1(n7976), .A2(n7827), .B1(n4172), .B2(n4890), .ZN(n1828)
         );
  AOI22_X1 U8308 ( .A1(n7977), .A2(n7827), .B1(n4692), .B2(n4892), .ZN(n1827)
         );
  AOI22_X1 U8309 ( .A1(n7978), .A2(n7827), .B1(n4173), .B2(n4894), .ZN(n1826)
         );
  AOI22_X1 U8310 ( .A1(n7979), .A2(n7827), .B1(n4693), .B2(n4896), .ZN(n1825)
         );
  AOI22_X1 U8311 ( .A1(n7980), .A2(n7827), .B1(n4382), .B2(n4898), .ZN(n1824)
         );
  AOI22_X1 U8312 ( .A1(n7981), .A2(n4844), .B1(n4383), .B2(n4900), .ZN(n1823)
         );
  AOI22_X1 U8313 ( .A1(n7982), .A2(n4844), .B1(n4694), .B2(n4902), .ZN(n1822)
         );
  AOI22_X1 U8314 ( .A1(n7983), .A2(n4844), .B1(n4174), .B2(n4904), .ZN(n1821)
         );
  AOI22_X1 U8315 ( .A1(n7984), .A2(n4844), .B1(n4175), .B2(n4906), .ZN(n1820)
         );
  AOI22_X1 U8316 ( .A1(n7985), .A2(n4844), .B1(n4695), .B2(n4908), .ZN(n1819)
         );
  NOR2_X1 U8317 ( .A1(alu_b_q[31]), .A2(n3831), .ZN(n7938) );
  AOI21_X1 U8318 ( .B1(alu_b_q[31]), .B2(n3831), .A(n7938), .ZN(n7940) );
  INV_X1 U8319 ( .A(n7940), .ZN(n7834) );
  OAI21_X1 U8320 ( .B1(alu_b_q[30]), .B2(n3833), .A(n7828), .ZN(n7932) );
  OAI21_X1 U8321 ( .B1(n7829), .B2(n7932), .A(n7933), .ZN(n7939) );
  XOR2_X1 U8322 ( .A(n7834), .B(n7939), .Z(n7862) );
  OAI22_X1 U8323 ( .A1(n3831), .A2(n7867), .B1(n7831), .B2(n7830), .ZN(n7832)
         );
  AOI211_X1 U8324 ( .C1(n7835), .C2(n7834), .A(n7833), .B(n7832), .ZN(n7850)
         );
  NOR4_X1 U8325 ( .A1(n7839), .A2(n7838), .A3(n7837), .A4(n7836), .ZN(n7841)
         );
  OAI22_X1 U8326 ( .A1(n7842), .A2(n7877), .B1(n7841), .B2(n7840), .ZN(n7848)
         );
  OAI22_X1 U8327 ( .A1(n7845), .A2(n7879), .B1(n7844), .B2(n7843), .ZN(n7847)
         );
  OAI21_X1 U8328 ( .B1(n7848), .B2(n7847), .A(n7846), .ZN(n7849) );
  OAI211_X1 U8329 ( .C1(n7852), .C2(n7851), .A(n7850), .B(n7849), .ZN(n7861)
         );
  AOI222_X1 U8330 ( .A1(n7853), .A2(alu_a_q[30]), .B1(n7853), .B2(alu_b_q[30]), 
        .C1(alu_a_q[30]), .C2(alu_b_q[30]), .ZN(n7854) );
  XOR2_X1 U8331 ( .A(n7854), .B(alu_a_q[31]), .Z(n7855) );
  XOR2_X1 U8332 ( .A(alu_b_q[31]), .B(n7855), .Z(n7859) );
  AOI21_X1 U8333 ( .B1(n7857), .B2(n7856), .A(n7872), .ZN(n7858) );
  OAI22_X1 U8334 ( .A1(n3842), .A2(n7859), .B1(n3873), .B2(n7858), .ZN(n7860)
         );
  AOI22_X1 U8335 ( .A1(n4847), .A2(n4845), .B1(n4696), .B2(n4846), .ZN(n1818)
         );
  AOI22_X1 U8336 ( .A1(n4849), .A2(n4845), .B1(n4384), .B2(n4848), .ZN(n1817)
         );
  AOI22_X1 U8337 ( .A1(n4851), .A2(n4845), .B1(n4385), .B2(n4850), .ZN(n1816)
         );
  AOI22_X1 U8338 ( .A1(n4853), .A2(n4845), .B1(n4386), .B2(n4852), .ZN(n1815)
         );
  AOI22_X1 U8339 ( .A1(n4855), .A2(n4845), .B1(n4700), .B2(n4854), .ZN(n1814)
         );
  AOI22_X1 U8340 ( .A1(n4857), .A2(n4845), .B1(n4176), .B2(n4856), .ZN(n1813)
         );
  AOI22_X1 U8341 ( .A1(n4859), .A2(n4845), .B1(n4177), .B2(n4858), .ZN(n1812)
         );
  AOI22_X1 U8342 ( .A1(n4861), .A2(n4845), .B1(n4701), .B2(n4860), .ZN(n1811)
         );
  AOI22_X1 U8343 ( .A1(n4863), .A2(n4845), .B1(n4697), .B2(n4862), .ZN(n1810)
         );
  AOI22_X1 U8344 ( .A1(n4865), .A2(n4845), .B1(n4387), .B2(n4864), .ZN(n1809)
         );
  AOI22_X1 U8345 ( .A1(n4867), .A2(n4845), .B1(n4388), .B2(n4866), .ZN(n1808)
         );
  AOI22_X1 U8346 ( .A1(n4869), .A2(n4845), .B1(n4389), .B2(n4868), .ZN(n1807)
         );
  AOI22_X1 U8347 ( .A1(n4871), .A2(n4845), .B1(n4702), .B2(n4870), .ZN(n1806)
         );
  AOI22_X1 U8348 ( .A1(n4873), .A2(n4845), .B1(n4178), .B2(n4872), .ZN(n1805)
         );
  AOI22_X1 U8349 ( .A1(n4875), .A2(n4845), .B1(n4179), .B2(n4874), .ZN(n1804)
         );
  AOI22_X1 U8350 ( .A1(n4877), .A2(n4845), .B1(n4703), .B2(n4876), .ZN(n1803)
         );
  AOI22_X1 U8351 ( .A1(n4879), .A2(n4845), .B1(n4698), .B2(n4878), .ZN(n1802)
         );
  AOI22_X1 U8352 ( .A1(n4881), .A2(n4845), .B1(n4390), .B2(n4880), .ZN(n1801)
         );
  AOI22_X1 U8353 ( .A1(n4883), .A2(n4845), .B1(n4391), .B2(n4882), .ZN(n1800)
         );
  AOI22_X1 U8354 ( .A1(n4885), .A2(n4845), .B1(n4392), .B2(n4884), .ZN(n1799)
         );
  AOI22_X1 U8355 ( .A1(n4887), .A2(n4845), .B1(n4704), .B2(n4886), .ZN(n1798)
         );
  AOI22_X1 U8356 ( .A1(n4889), .A2(n7863), .B1(n4180), .B2(n4888), .ZN(n1797)
         );
  AOI22_X1 U8357 ( .A1(n4891), .A2(n7863), .B1(n4181), .B2(n4890), .ZN(n1796)
         );
  AOI22_X1 U8358 ( .A1(n4893), .A2(n7863), .B1(n4705), .B2(n4892), .ZN(n1795)
         );
  AOI22_X1 U8359 ( .A1(n4895), .A2(n7863), .B1(n4699), .B2(n4894), .ZN(n1794)
         );
  AOI22_X1 U8360 ( .A1(n4897), .A2(n7863), .B1(n4393), .B2(n4896), .ZN(n1793)
         );
  AOI22_X1 U8361 ( .A1(n4899), .A2(n7863), .B1(n4394), .B2(n4898), .ZN(n1792)
         );
  AOI22_X1 U8362 ( .A1(n4901), .A2(n4845), .B1(n4395), .B2(n4900), .ZN(n1791)
         );
  AOI22_X1 U8363 ( .A1(n4903), .A2(n4845), .B1(n4706), .B2(n4902), .ZN(n1790)
         );
  AOI22_X1 U8364 ( .A1(n4905), .A2(n4845), .B1(n4182), .B2(n4904), .ZN(n1789)
         );
  AOI22_X1 U8365 ( .A1(n4907), .A2(n4845), .B1(n4183), .B2(n4906), .ZN(n1788)
         );
  AOI22_X1 U8366 ( .A1(n4909), .A2(n4845), .B1(n4707), .B2(n4908), .ZN(n1787)
         );
  NAND2_X1 U8367 ( .A1(n7865), .A2(n7864), .ZN(n7875) );
  INV_X1 U8368 ( .A(n7875), .ZN(n7869) );
  OAI21_X1 U8369 ( .B1(n7866), .B2(n7885), .A(n3807), .ZN(n7868) );
  OAI221_X1 U8370 ( .B1(alu_b_q[0]), .B2(n7869), .C1(alu_b_q[0]), .C2(n7868), 
        .A(n7867), .ZN(n7953) );
  AOI22_X1 U8371 ( .A1(alu_b_q[0]), .A2(n7872), .B1(n7871), .B2(n7870), .ZN(
        n7951) );
  AOI22_X1 U8372 ( .A1(n7876), .A2(n7875), .B1(n7874), .B2(n7873), .ZN(n7950)
         );
  OAI22_X1 U8373 ( .A1(n7880), .A2(n7879), .B1(n7878), .B2(n7877), .ZN(n7886)
         );
  OAI211_X1 U8374 ( .C1(n7883), .C2(n3803), .A(n7882), .B(n7881), .ZN(n7884)
         );
  AOI22_X1 U8375 ( .A1(n7887), .A2(n7886), .B1(n7885), .B2(n7884), .ZN(n7949)
         );
  NOR4_X1 U8376 ( .A1(n7938), .A2(n7889), .A3(n7888), .A4(n7932), .ZN(n7937)
         );
  NAND2_X1 U8377 ( .A1(alu_b_q[20]), .A2(n3791), .ZN(n7920) );
  NOR2_X1 U8378 ( .A1(n7891), .A2(n7890), .ZN(n7913) );
  NOR2_X1 U8379 ( .A1(alu_a_q[11]), .A2(n3775), .ZN(n7894) );
  OAI21_X1 U8380 ( .B1(n7894), .B2(n7893), .A(n7892), .ZN(n7898) );
  OR2_X1 U8381 ( .A1(n7905), .A2(n7895), .ZN(n7896) );
  AOI221_X1 U8382 ( .B1(n7899), .B2(n7898), .C1(n7897), .C2(n7898), .A(n7896), 
        .ZN(n7909) );
  NOR2_X1 U8383 ( .A1(alu_a_q[13]), .A2(n3776), .ZN(n7900) );
  AOI211_X1 U8384 ( .C1(n7903), .C2(n7902), .A(n7901), .B(n7900), .ZN(n7906)
         );
  OAI21_X1 U8385 ( .B1(n7906), .B2(n7905), .A(n7904), .ZN(n7908) );
  OAI21_X1 U8386 ( .B1(n7909), .B2(n7908), .A(n7907), .ZN(n7912) );
  OAI21_X1 U8387 ( .B1(alu_b_q[18]), .B2(n3786), .A(n7910), .ZN(n7911) );
  AOI21_X1 U8388 ( .B1(n7913), .B2(n7912), .A(n7911), .ZN(n7916) );
  OAI211_X1 U8389 ( .C1(n7917), .C2(n7916), .A(n7915), .B(n7914), .ZN(n7919)
         );
  OAI221_X1 U8390 ( .B1(n7921), .B2(n7920), .C1(n7921), .C2(n7919), .A(n7918), 
        .ZN(n7922) );
  OAI211_X1 U8391 ( .C1(alu_b_q[22]), .C2(n3795), .A(n7923), .B(n7922), .ZN(
        n7925) );
  NAND2_X1 U8392 ( .A1(alu_b_q[25]), .A2(n3829), .ZN(n7924) );
  OAI221_X1 U8393 ( .B1(n7927), .B2(n7926), .C1(n7927), .C2(n7925), .A(n7924), 
        .ZN(n7936) );
  AOI211_X1 U8394 ( .C1(n7931), .C2(n7930), .A(n7929), .B(n7928), .ZN(n7934)
         );
  AOI221_X1 U8395 ( .B1(n7934), .B2(n7933), .C1(n7932), .C2(n7933), .A(n7938), 
        .ZN(n7935) );
  AOI211_X1 U8396 ( .C1(n7937), .C2(n7936), .A(n7935), .B(n3830), .ZN(n7944)
         );
  NAND2_X1 U8397 ( .A1(alu_b_q[31]), .A2(n3831), .ZN(n7943) );
  AOI211_X1 U8398 ( .C1(n7940), .C2(n7939), .A(n157), .B(n7938), .ZN(n7942) );
  AOI211_X1 U8399 ( .C1(n7944), .C2(n7943), .A(n7942), .B(n7941), .ZN(n7945)
         );
  AOI22_X1 U8400 ( .A1(n7947), .A2(n7946), .B1(n7945), .B2(n3835), .ZN(n7948)
         );
  NAND4_X1 U8401 ( .A1(n7951), .A2(n7950), .A3(n7949), .A4(n7948), .ZN(n7952)
         );
endmodule

